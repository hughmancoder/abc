// Benchmark "adder" written by ABC on Sun Jun 22 16:29:23 2025

module adder ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n387, new_n388, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n413, new_n414, new_n415, new_n416, new_n417, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n427,
    new_n428, new_n429, new_n430, new_n431, new_n432, new_n433, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n451,
    new_n452, new_n453, new_n454, new_n455, new_n456, new_n457, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n483,
    new_n484, new_n485, new_n486, new_n487, new_n488, new_n489, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1323, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1371, new_n1372,
    new_n1373, new_n1374, new_n1375, new_n1376, new_n1377, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1387, new_n1388, new_n1389, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1515, new_n1516, new_n1517, new_n1518,
    new_n1519, new_n1520, new_n1521, new_n1522, new_n1523, new_n1524,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1532, new_n1533, new_n1534, new_n1535, new_n1536,
    new_n1537, new_n1538, new_n1539, new_n1540, new_n1541, new_n1542,
    new_n1543, new_n1544, new_n1545, new_n1546, new_n1547, new_n1548,
    new_n1549, new_n1550, new_n1551, new_n1552, new_n1553, new_n1554,
    new_n1555, new_n1556, new_n1557, new_n1558, new_n1559, new_n1560,
    new_n1561, new_n1562, new_n1563, new_n1564, new_n1565, new_n1566,
    new_n1567, new_n1568, new_n1569, new_n1570, new_n1571, new_n1572,
    new_n1573, new_n1574, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1584, new_n1585,
    new_n1586;
  XOR2_HPNW1   g0000(.A(\b[0] ), .B(\a[0] ), .Y(\f[0] ));
  INV1_HPNW1   g0001(.A(\b[1] ), .Y(new_n387));
  NAND2_HPNW1  g0002(.A(\b[0] ), .B(\a[0] ), .Y(new_n388));
  XOR3_HPNW1   g0003(.A(new_n388), .B(new_n387), .C(\a[1] ), .Y(\f[1] ));
  AND2_HPNW1   g0004(.A(\b[1] ), .B(\a[1] ), .Y(new_n390));
  NOR2_HPNW1   g0005(.A(\b[1] ), .B(\a[1] ), .Y(new_n391));
  NOR2_HPNW1   g0006(.A(new_n391), .B(new_n388), .Y(new_n392));
  NOR2_HPNW1   g0007(.A(new_n390), .B(new_n392), .Y(new_n393));
  OR2_HPNW1    g0008(.A(\a[2] ), .B(\b[2] ), .Y(new_n394));
  NAND2_HPNW1  g0009(.A(\b[2] ), .B(\a[2] ), .Y(new_n395));
  NAND2_HPNW1  g0010(.A(new_n394), .B(new_n395), .Y(new_n396));
  XOR2_HPNW1   g0011(.A(new_n396), .B(new_n393), .Y(\f[2] ));
  INV1_HPNW1   g0012(.A(new_n394), .Y(new_n398));
  OAI21_HPNW1  g0013(.A0(new_n398), .A1(new_n393), .B0(new_n395), .Y(new_n399));
  INV1_HPNW1   g0014(.A(\a[3] ), .Y(new_n400));
  INV1_HPNW1   g0015(.A(\b[3] ), .Y(new_n401));
  NAND2_HPNW1  g0016(.A(new_n401), .B(new_n400), .Y(new_n402));
  NAND2_HPNW1  g0017(.A(\b[3] ), .B(\a[3] ), .Y(new_n403));
  NAND2_HPNW1  g0018(.A(new_n402), .B(new_n403), .Y(new_n404));
  XNOR2_HPNW1  g0019(.A(new_n399), .B(new_n404), .Y(\f[3] ));
  INV1_HPNW1   g0020(.A(new_n403), .Y(new_n406));
  AOI21_HPNW1  g0021(.A0(new_n402), .A1(new_n399), .B0(new_n406), .Y(new_n407));
  NOR2_HPNW1   g0022(.A(\b[4] ), .B(\a[4] ), .Y(new_n408));
  INV1_HPNW1   g0023(.A(new_n408), .Y(new_n409));
  NAND2_HPNW1  g0024(.A(\b[4] ), .B(\a[4] ), .Y(new_n410));
  NAND2_HPNW1  g0025(.A(new_n409), .B(new_n410), .Y(new_n411));
  XOR2_HPNW1   g0026(.A(new_n411), .B(new_n407), .Y(\f[4] ));
  OAI21_HPNW1  g0027(.A0(new_n408), .A1(new_n407), .B0(new_n410), .Y(new_n413));
  NOR2_HPNW1   g0028(.A(\b[5] ), .B(\a[5] ), .Y(new_n414));
  INV1_HPNW1   g0029(.A(new_n414), .Y(new_n415));
  NAND2_HPNW1  g0030(.A(\b[5] ), .B(\a[5] ), .Y(new_n416));
  NAND2_HPNW1  g0031(.A(new_n415), .B(new_n416), .Y(new_n417));
  XNOR2_HPNW1  g0032(.A(new_n413), .B(new_n417), .Y(\f[5] ));
  INV1_HPNW1   g0033(.A(new_n416), .Y(new_n419));
  AOI21_HPNW1  g0034(.A0(new_n415), .A1(new_n413), .B0(new_n419), .Y(new_n420));
  INV1_HPNW1   g0035(.A(\a[6] ), .Y(new_n421));
  INV1_HPNW1   g0036(.A(\b[6] ), .Y(new_n422));
  NAND2_HPNW1  g0037(.A(new_n422), .B(new_n421), .Y(new_n423));
  NAND2_HPNW1  g0038(.A(\b[6] ), .B(\a[6] ), .Y(new_n424));
  NAND2_HPNW1  g0039(.A(new_n423), .B(new_n424), .Y(new_n425));
  XOR2_HPNW1   g0040(.A(new_n425), .B(new_n420), .Y(\f[6] ));
  INV1_HPNW1   g0041(.A(new_n423), .Y(new_n427));
  OAI21_HPNW1  g0042(.A0(new_n427), .A1(new_n420), .B0(new_n424), .Y(new_n428));
  INV1_HPNW1   g0043(.A(\a[7] ), .Y(new_n429));
  INV1_HPNW1   g0044(.A(\b[7] ), .Y(new_n430));
  NAND2_HPNW1  g0045(.A(new_n430), .B(new_n429), .Y(new_n431));
  NAND2_HPNW1  g0046(.A(\b[7] ), .B(\a[7] ), .Y(new_n432));
  NAND2_HPNW1  g0047(.A(new_n431), .B(new_n432), .Y(new_n433));
  XNOR2_HPNW1  g0048(.A(new_n428), .B(new_n433), .Y(\f[7] ));
  INV1_HPNW1   g0049(.A(new_n432), .Y(new_n435));
  AOI21_HPNW1  g0050(.A0(new_n431), .A1(new_n428), .B0(new_n435), .Y(new_n436));
  INV1_HPNW1   g0051(.A(\a[8] ), .Y(new_n437));
  INV1_HPNW1   g0052(.A(\b[8] ), .Y(new_n438));
  NAND2_HPNW1  g0053(.A(new_n438), .B(new_n437), .Y(new_n439));
  NAND2_HPNW1  g0054(.A(\b[8] ), .B(\a[8] ), .Y(new_n440));
  NAND2_HPNW1  g0055(.A(new_n439), .B(new_n440), .Y(new_n441));
  XOR2_HPNW1   g0056(.A(new_n441), .B(new_n436), .Y(\f[8] ));
  INV1_HPNW1   g0057(.A(new_n439), .Y(new_n443));
  OAI21_HPNW1  g0058(.A0(new_n443), .A1(new_n436), .B0(new_n440), .Y(new_n444));
  INV1_HPNW1   g0059(.A(\a[9] ), .Y(new_n445));
  INV1_HPNW1   g0060(.A(\b[9] ), .Y(new_n446));
  NAND2_HPNW1  g0061(.A(new_n446), .B(new_n445), .Y(new_n447));
  NAND2_HPNW1  g0062(.A(\b[9] ), .B(\a[9] ), .Y(new_n448));
  NAND2_HPNW1  g0063(.A(new_n447), .B(new_n448), .Y(new_n449));
  XNOR2_HPNW1  g0064(.A(new_n444), .B(new_n449), .Y(\f[9] ));
  INV1_HPNW1   g0065(.A(new_n448), .Y(new_n451));
  AOI21_HPNW1  g0066(.A0(new_n447), .A1(new_n444), .B0(new_n451), .Y(new_n452));
  INV1_HPNW1   g0067(.A(\a[10] ), .Y(new_n453));
  INV1_HPNW1   g0068(.A(\b[10] ), .Y(new_n454));
  NAND2_HPNW1  g0069(.A(new_n454), .B(new_n453), .Y(new_n455));
  NAND2_HPNW1  g0070(.A(\b[10] ), .B(\a[10] ), .Y(new_n456));
  NAND2_HPNW1  g0071(.A(new_n455), .B(new_n456), .Y(new_n457));
  XOR2_HPNW1   g0072(.A(new_n457), .B(new_n452), .Y(\f[10] ));
  INV1_HPNW1   g0073(.A(new_n455), .Y(new_n459));
  OAI21_HPNW1  g0074(.A0(new_n459), .A1(new_n452), .B0(new_n456), .Y(new_n460));
  INV1_HPNW1   g0075(.A(\a[11] ), .Y(new_n461));
  INV1_HPNW1   g0076(.A(\b[11] ), .Y(new_n462));
  NAND2_HPNW1  g0077(.A(new_n462), .B(new_n461), .Y(new_n463));
  NAND2_HPNW1  g0078(.A(\b[11] ), .B(\a[11] ), .Y(new_n464));
  NAND2_HPNW1  g0079(.A(new_n463), .B(new_n464), .Y(new_n465));
  XNOR2_HPNW1  g0080(.A(new_n460), .B(new_n465), .Y(\f[11] ));
  INV1_HPNW1   g0081(.A(new_n464), .Y(new_n467));
  AOI21_HPNW1  g0082(.A0(new_n463), .A1(new_n460), .B0(new_n467), .Y(new_n468));
  INV1_HPNW1   g0083(.A(\a[12] ), .Y(new_n469));
  INV1_HPNW1   g0084(.A(\b[12] ), .Y(new_n470));
  NAND2_HPNW1  g0085(.A(new_n470), .B(new_n469), .Y(new_n471));
  NAND2_HPNW1  g0086(.A(\b[12] ), .B(\a[12] ), .Y(new_n472));
  NAND2_HPNW1  g0087(.A(new_n471), .B(new_n472), .Y(new_n473));
  XOR2_HPNW1   g0088(.A(new_n473), .B(new_n468), .Y(\f[12] ));
  INV1_HPNW1   g0089(.A(new_n471), .Y(new_n475));
  OAI21_HPNW1  g0090(.A0(new_n475), .A1(new_n468), .B0(new_n472), .Y(new_n476));
  INV1_HPNW1   g0091(.A(\a[13] ), .Y(new_n477));
  INV1_HPNW1   g0092(.A(\b[13] ), .Y(new_n478));
  NAND2_HPNW1  g0093(.A(new_n478), .B(new_n477), .Y(new_n479));
  NAND2_HPNW1  g0094(.A(\b[13] ), .B(\a[13] ), .Y(new_n480));
  NAND2_HPNW1  g0095(.A(new_n479), .B(new_n480), .Y(new_n481));
  XNOR2_HPNW1  g0096(.A(new_n476), .B(new_n481), .Y(\f[13] ));
  INV1_HPNW1   g0097(.A(new_n480), .Y(new_n483));
  AOI21_HPNW1  g0098(.A0(new_n479), .A1(new_n476), .B0(new_n483), .Y(new_n484));
  INV1_HPNW1   g0099(.A(\a[14] ), .Y(new_n485));
  INV1_HPNW1   g0100(.A(\b[14] ), .Y(new_n486));
  NAND2_HPNW1  g0101(.A(new_n486), .B(new_n485), .Y(new_n487));
  NAND2_HPNW1  g0102(.A(\b[14] ), .B(\a[14] ), .Y(new_n488));
  NAND2_HPNW1  g0103(.A(new_n487), .B(new_n488), .Y(new_n489));
  XOR2_HPNW1   g0104(.A(new_n489), .B(new_n484), .Y(\f[14] ));
  INV1_HPNW1   g0105(.A(new_n487), .Y(new_n491));
  OAI21_HPNW1  g0106(.A0(new_n491), .A1(new_n484), .B0(new_n488), .Y(new_n492));
  INV1_HPNW1   g0107(.A(\a[15] ), .Y(new_n493));
  INV1_HPNW1   g0108(.A(\b[15] ), .Y(new_n494));
  NAND2_HPNW1  g0109(.A(new_n494), .B(new_n493), .Y(new_n495));
  NAND2_HPNW1  g0110(.A(\b[15] ), .B(\a[15] ), .Y(new_n496));
  NAND2_HPNW1  g0111(.A(new_n495), .B(new_n496), .Y(new_n497));
  XNOR2_HPNW1  g0112(.A(new_n492), .B(new_n497), .Y(\f[15] ));
  INV1_HPNW1   g0113(.A(new_n496), .Y(new_n499));
  AOI21_HPNW1  g0114(.A0(new_n495), .A1(new_n492), .B0(new_n499), .Y(new_n500));
  INV1_HPNW1   g0115(.A(\a[16] ), .Y(new_n501));
  INV1_HPNW1   g0116(.A(\b[16] ), .Y(new_n502));
  NAND2_HPNW1  g0117(.A(new_n502), .B(new_n501), .Y(new_n503));
  NAND2_HPNW1  g0118(.A(\b[16] ), .B(\a[16] ), .Y(new_n504));
  NAND2_HPNW1  g0119(.A(new_n503), .B(new_n504), .Y(new_n505));
  XOR2_HPNW1   g0120(.A(new_n505), .B(new_n500), .Y(\f[16] ));
  INV1_HPNW1   g0121(.A(new_n503), .Y(new_n507));
  OAI21_HPNW1  g0122(.A0(new_n507), .A1(new_n500), .B0(new_n504), .Y(new_n508));
  INV1_HPNW1   g0123(.A(\a[17] ), .Y(new_n509));
  INV1_HPNW1   g0124(.A(\b[17] ), .Y(new_n510));
  NAND2_HPNW1  g0125(.A(new_n510), .B(new_n509), .Y(new_n511));
  NAND2_HPNW1  g0126(.A(\b[17] ), .B(\a[17] ), .Y(new_n512));
  NAND2_HPNW1  g0127(.A(new_n511), .B(new_n512), .Y(new_n513));
  XNOR2_HPNW1  g0128(.A(new_n508), .B(new_n513), .Y(\f[17] ));
  INV1_HPNW1   g0129(.A(new_n512), .Y(new_n515));
  AOI21_HPNW1  g0130(.A0(new_n511), .A1(new_n508), .B0(new_n515), .Y(new_n516));
  INV1_HPNW1   g0131(.A(\a[18] ), .Y(new_n517));
  INV1_HPNW1   g0132(.A(\b[18] ), .Y(new_n518));
  NAND2_HPNW1  g0133(.A(new_n518), .B(new_n517), .Y(new_n519));
  NAND2_HPNW1  g0134(.A(\b[18] ), .B(\a[18] ), .Y(new_n520));
  NAND2_HPNW1  g0135(.A(new_n519), .B(new_n520), .Y(new_n521));
  XOR2_HPNW1   g0136(.A(new_n521), .B(new_n516), .Y(\f[18] ));
  INV1_HPNW1   g0137(.A(new_n519), .Y(new_n523));
  OAI21_HPNW1  g0138(.A0(new_n523), .A1(new_n516), .B0(new_n520), .Y(new_n524));
  INV1_HPNW1   g0139(.A(\a[19] ), .Y(new_n525));
  INV1_HPNW1   g0140(.A(\b[19] ), .Y(new_n526));
  NAND2_HPNW1  g0141(.A(new_n526), .B(new_n525), .Y(new_n527));
  NAND2_HPNW1  g0142(.A(\b[19] ), .B(\a[19] ), .Y(new_n528));
  NAND2_HPNW1  g0143(.A(new_n527), .B(new_n528), .Y(new_n529));
  XNOR2_HPNW1  g0144(.A(new_n524), .B(new_n529), .Y(\f[19] ));
  INV1_HPNW1   g0145(.A(new_n528), .Y(new_n531));
  AOI21_HPNW1  g0146(.A0(new_n527), .A1(new_n524), .B0(new_n531), .Y(new_n532));
  INV1_HPNW1   g0147(.A(\a[20] ), .Y(new_n533));
  INV1_HPNW1   g0148(.A(\b[20] ), .Y(new_n534));
  NAND2_HPNW1  g0149(.A(new_n534), .B(new_n533), .Y(new_n535));
  NAND2_HPNW1  g0150(.A(\b[20] ), .B(\a[20] ), .Y(new_n536));
  NAND2_HPNW1  g0151(.A(new_n535), .B(new_n536), .Y(new_n537));
  XOR2_HPNW1   g0152(.A(new_n537), .B(new_n532), .Y(\f[20] ));
  INV1_HPNW1   g0153(.A(new_n535), .Y(new_n539));
  OAI21_HPNW1  g0154(.A0(new_n539), .A1(new_n532), .B0(new_n536), .Y(new_n540));
  INV1_HPNW1   g0155(.A(\a[21] ), .Y(new_n541));
  INV1_HPNW1   g0156(.A(\b[21] ), .Y(new_n542));
  NAND2_HPNW1  g0157(.A(new_n542), .B(new_n541), .Y(new_n543));
  NAND2_HPNW1  g0158(.A(\b[21] ), .B(\a[21] ), .Y(new_n544));
  NAND2_HPNW1  g0159(.A(new_n543), .B(new_n544), .Y(new_n545));
  XNOR2_HPNW1  g0160(.A(new_n540), .B(new_n545), .Y(\f[21] ));
  INV1_HPNW1   g0161(.A(new_n544), .Y(new_n547));
  AOI21_HPNW1  g0162(.A0(new_n543), .A1(new_n540), .B0(new_n547), .Y(new_n548));
  INV1_HPNW1   g0163(.A(\a[22] ), .Y(new_n549));
  INV1_HPNW1   g0164(.A(\b[22] ), .Y(new_n550));
  NAND2_HPNW1  g0165(.A(new_n550), .B(new_n549), .Y(new_n551));
  NAND2_HPNW1  g0166(.A(\b[22] ), .B(\a[22] ), .Y(new_n552));
  NAND2_HPNW1  g0167(.A(new_n551), .B(new_n552), .Y(new_n553));
  XOR2_HPNW1   g0168(.A(new_n553), .B(new_n548), .Y(\f[22] ));
  INV1_HPNW1   g0169(.A(new_n551), .Y(new_n555));
  OAI21_HPNW1  g0170(.A0(new_n555), .A1(new_n548), .B0(new_n552), .Y(new_n556));
  INV1_HPNW1   g0171(.A(\a[23] ), .Y(new_n557));
  INV1_HPNW1   g0172(.A(\b[23] ), .Y(new_n558));
  NAND2_HPNW1  g0173(.A(new_n558), .B(new_n557), .Y(new_n559));
  NAND2_HPNW1  g0174(.A(\b[23] ), .B(\a[23] ), .Y(new_n560));
  NAND2_HPNW1  g0175(.A(new_n559), .B(new_n560), .Y(new_n561));
  XNOR2_HPNW1  g0176(.A(new_n556), .B(new_n561), .Y(\f[23] ));
  INV1_HPNW1   g0177(.A(new_n560), .Y(new_n563));
  AOI21_HPNW1  g0178(.A0(new_n559), .A1(new_n556), .B0(new_n563), .Y(new_n564));
  INV1_HPNW1   g0179(.A(\a[24] ), .Y(new_n565));
  INV1_HPNW1   g0180(.A(\b[24] ), .Y(new_n566));
  NAND2_HPNW1  g0181(.A(new_n566), .B(new_n565), .Y(new_n567));
  NAND2_HPNW1  g0182(.A(\b[24] ), .B(\a[24] ), .Y(new_n568));
  NAND2_HPNW1  g0183(.A(new_n567), .B(new_n568), .Y(new_n569));
  XOR2_HPNW1   g0184(.A(new_n569), .B(new_n564), .Y(\f[24] ));
  INV1_HPNW1   g0185(.A(new_n567), .Y(new_n571));
  OAI21_HPNW1  g0186(.A0(new_n571), .A1(new_n564), .B0(new_n568), .Y(new_n572));
  INV1_HPNW1   g0187(.A(\a[25] ), .Y(new_n573));
  INV1_HPNW1   g0188(.A(\b[25] ), .Y(new_n574));
  NAND2_HPNW1  g0189(.A(new_n574), .B(new_n573), .Y(new_n575));
  NAND2_HPNW1  g0190(.A(\b[25] ), .B(\a[25] ), .Y(new_n576));
  NAND2_HPNW1  g0191(.A(new_n575), .B(new_n576), .Y(new_n577));
  XNOR2_HPNW1  g0192(.A(new_n572), .B(new_n577), .Y(\f[25] ));
  INV1_HPNW1   g0193(.A(new_n576), .Y(new_n579));
  AOI21_HPNW1  g0194(.A0(new_n575), .A1(new_n572), .B0(new_n579), .Y(new_n580));
  INV1_HPNW1   g0195(.A(\a[26] ), .Y(new_n581));
  INV1_HPNW1   g0196(.A(\b[26] ), .Y(new_n582));
  NAND2_HPNW1  g0197(.A(new_n582), .B(new_n581), .Y(new_n583));
  NAND2_HPNW1  g0198(.A(\b[26] ), .B(\a[26] ), .Y(new_n584));
  NAND2_HPNW1  g0199(.A(new_n583), .B(new_n584), .Y(new_n585));
  XOR2_HPNW1   g0200(.A(new_n585), .B(new_n580), .Y(\f[26] ));
  INV1_HPNW1   g0201(.A(new_n583), .Y(new_n587));
  OAI21_HPNW1  g0202(.A0(new_n587), .A1(new_n580), .B0(new_n584), .Y(new_n588));
  INV1_HPNW1   g0203(.A(\a[27] ), .Y(new_n589));
  INV1_HPNW1   g0204(.A(\b[27] ), .Y(new_n590));
  NAND2_HPNW1  g0205(.A(new_n590), .B(new_n589), .Y(new_n591));
  NAND2_HPNW1  g0206(.A(\b[27] ), .B(\a[27] ), .Y(new_n592));
  NAND2_HPNW1  g0207(.A(new_n591), .B(new_n592), .Y(new_n593));
  XNOR2_HPNW1  g0208(.A(new_n588), .B(new_n593), .Y(\f[27] ));
  INV1_HPNW1   g0209(.A(new_n592), .Y(new_n595));
  AOI21_HPNW1  g0210(.A0(new_n591), .A1(new_n588), .B0(new_n595), .Y(new_n596));
  INV1_HPNW1   g0211(.A(\a[28] ), .Y(new_n597));
  INV1_HPNW1   g0212(.A(\b[28] ), .Y(new_n598));
  NAND2_HPNW1  g0213(.A(new_n598), .B(new_n597), .Y(new_n599));
  NAND2_HPNW1  g0214(.A(\b[28] ), .B(\a[28] ), .Y(new_n600));
  NAND2_HPNW1  g0215(.A(new_n599), .B(new_n600), .Y(new_n601));
  XOR2_HPNW1   g0216(.A(new_n601), .B(new_n596), .Y(\f[28] ));
  INV1_HPNW1   g0217(.A(new_n599), .Y(new_n603));
  OAI21_HPNW1  g0218(.A0(new_n603), .A1(new_n596), .B0(new_n600), .Y(new_n604));
  INV1_HPNW1   g0219(.A(\a[29] ), .Y(new_n605));
  INV1_HPNW1   g0220(.A(\b[29] ), .Y(new_n606));
  NAND2_HPNW1  g0221(.A(new_n606), .B(new_n605), .Y(new_n607));
  NAND2_HPNW1  g0222(.A(\b[29] ), .B(\a[29] ), .Y(new_n608));
  NAND2_HPNW1  g0223(.A(new_n607), .B(new_n608), .Y(new_n609));
  XNOR2_HPNW1  g0224(.A(new_n604), .B(new_n609), .Y(\f[29] ));
  INV1_HPNW1   g0225(.A(new_n608), .Y(new_n611));
  AOI21_HPNW1  g0226(.A0(new_n607), .A1(new_n604), .B0(new_n611), .Y(new_n612));
  INV1_HPNW1   g0227(.A(\a[30] ), .Y(new_n613));
  INV1_HPNW1   g0228(.A(\b[30] ), .Y(new_n614));
  NAND2_HPNW1  g0229(.A(new_n614), .B(new_n613), .Y(new_n615));
  NAND2_HPNW1  g0230(.A(\b[30] ), .B(\a[30] ), .Y(new_n616));
  NAND2_HPNW1  g0231(.A(new_n615), .B(new_n616), .Y(new_n617));
  XOR2_HPNW1   g0232(.A(new_n617), .B(new_n612), .Y(\f[30] ));
  INV1_HPNW1   g0233(.A(new_n615), .Y(new_n619));
  OAI21_HPNW1  g0234(.A0(new_n619), .A1(new_n612), .B0(new_n616), .Y(new_n620));
  INV1_HPNW1   g0235(.A(\a[31] ), .Y(new_n621));
  INV1_HPNW1   g0236(.A(\b[31] ), .Y(new_n622));
  NAND2_HPNW1  g0237(.A(new_n622), .B(new_n621), .Y(new_n623));
  NAND2_HPNW1  g0238(.A(\b[31] ), .B(\a[31] ), .Y(new_n624));
  NAND2_HPNW1  g0239(.A(new_n623), .B(new_n624), .Y(new_n625));
  XNOR2_HPNW1  g0240(.A(new_n620), .B(new_n625), .Y(\f[31] ));
  INV1_HPNW1   g0241(.A(new_n624), .Y(new_n627));
  AOI21_HPNW1  g0242(.A0(new_n623), .A1(new_n620), .B0(new_n627), .Y(new_n628));
  INV1_HPNW1   g0243(.A(\a[32] ), .Y(new_n629));
  INV1_HPNW1   g0244(.A(\b[32] ), .Y(new_n630));
  NAND2_HPNW1  g0245(.A(new_n630), .B(new_n629), .Y(new_n631));
  NAND2_HPNW1  g0246(.A(\b[32] ), .B(\a[32] ), .Y(new_n632));
  NAND2_HPNW1  g0247(.A(new_n631), .B(new_n632), .Y(new_n633));
  XOR2_HPNW1   g0248(.A(new_n633), .B(new_n628), .Y(\f[32] ));
  INV1_HPNW1   g0249(.A(new_n631), .Y(new_n635));
  OAI21_HPNW1  g0250(.A0(new_n635), .A1(new_n628), .B0(new_n632), .Y(new_n636));
  INV1_HPNW1   g0251(.A(\a[33] ), .Y(new_n637));
  INV1_HPNW1   g0252(.A(\b[33] ), .Y(new_n638));
  NAND2_HPNW1  g0253(.A(new_n638), .B(new_n637), .Y(new_n639));
  NAND2_HPNW1  g0254(.A(\b[33] ), .B(\a[33] ), .Y(new_n640));
  NAND2_HPNW1  g0255(.A(new_n639), .B(new_n640), .Y(new_n641));
  XNOR2_HPNW1  g0256(.A(new_n636), .B(new_n641), .Y(\f[33] ));
  INV1_HPNW1   g0257(.A(new_n640), .Y(new_n643));
  AOI21_HPNW1  g0258(.A0(new_n639), .A1(new_n636), .B0(new_n643), .Y(new_n644));
  INV1_HPNW1   g0259(.A(\a[34] ), .Y(new_n645));
  INV1_HPNW1   g0260(.A(\b[34] ), .Y(new_n646));
  NAND2_HPNW1  g0261(.A(new_n646), .B(new_n645), .Y(new_n647));
  NAND2_HPNW1  g0262(.A(\b[34] ), .B(\a[34] ), .Y(new_n648));
  NAND2_HPNW1  g0263(.A(new_n647), .B(new_n648), .Y(new_n649));
  XOR2_HPNW1   g0264(.A(new_n649), .B(new_n644), .Y(\f[34] ));
  INV1_HPNW1   g0265(.A(new_n647), .Y(new_n651));
  OAI21_HPNW1  g0266(.A0(new_n651), .A1(new_n644), .B0(new_n648), .Y(new_n652));
  INV1_HPNW1   g0267(.A(\a[35] ), .Y(new_n653));
  INV1_HPNW1   g0268(.A(\b[35] ), .Y(new_n654));
  NAND2_HPNW1  g0269(.A(new_n654), .B(new_n653), .Y(new_n655));
  NAND2_HPNW1  g0270(.A(\b[35] ), .B(\a[35] ), .Y(new_n656));
  NAND2_HPNW1  g0271(.A(new_n655), .B(new_n656), .Y(new_n657));
  XNOR2_HPNW1  g0272(.A(new_n652), .B(new_n657), .Y(\f[35] ));
  INV1_HPNW1   g0273(.A(new_n656), .Y(new_n659));
  AOI21_HPNW1  g0274(.A0(new_n655), .A1(new_n652), .B0(new_n659), .Y(new_n660));
  INV1_HPNW1   g0275(.A(\a[36] ), .Y(new_n661));
  INV1_HPNW1   g0276(.A(\b[36] ), .Y(new_n662));
  NAND2_HPNW1  g0277(.A(new_n662), .B(new_n661), .Y(new_n663));
  NAND2_HPNW1  g0278(.A(\b[36] ), .B(\a[36] ), .Y(new_n664));
  NAND2_HPNW1  g0279(.A(new_n663), .B(new_n664), .Y(new_n665));
  XOR2_HPNW1   g0280(.A(new_n665), .B(new_n660), .Y(\f[36] ));
  INV1_HPNW1   g0281(.A(new_n663), .Y(new_n667));
  OAI21_HPNW1  g0282(.A0(new_n667), .A1(new_n660), .B0(new_n664), .Y(new_n668));
  INV1_HPNW1   g0283(.A(\a[37] ), .Y(new_n669));
  INV1_HPNW1   g0284(.A(\b[37] ), .Y(new_n670));
  NAND2_HPNW1  g0285(.A(new_n670), .B(new_n669), .Y(new_n671));
  NAND2_HPNW1  g0286(.A(\b[37] ), .B(\a[37] ), .Y(new_n672));
  NAND2_HPNW1  g0287(.A(new_n671), .B(new_n672), .Y(new_n673));
  XNOR2_HPNW1  g0288(.A(new_n668), .B(new_n673), .Y(\f[37] ));
  INV1_HPNW1   g0289(.A(new_n672), .Y(new_n675));
  AOI21_HPNW1  g0290(.A0(new_n671), .A1(new_n668), .B0(new_n675), .Y(new_n676));
  INV1_HPNW1   g0291(.A(\a[38] ), .Y(new_n677));
  INV1_HPNW1   g0292(.A(\b[38] ), .Y(new_n678));
  NAND2_HPNW1  g0293(.A(new_n678), .B(new_n677), .Y(new_n679));
  NAND2_HPNW1  g0294(.A(\b[38] ), .B(\a[38] ), .Y(new_n680));
  NAND2_HPNW1  g0295(.A(new_n679), .B(new_n680), .Y(new_n681));
  XOR2_HPNW1   g0296(.A(new_n681), .B(new_n676), .Y(\f[38] ));
  INV1_HPNW1   g0297(.A(new_n679), .Y(new_n683));
  OAI21_HPNW1  g0298(.A0(new_n683), .A1(new_n676), .B0(new_n680), .Y(new_n684));
  INV1_HPNW1   g0299(.A(\a[39] ), .Y(new_n685));
  INV1_HPNW1   g0300(.A(\b[39] ), .Y(new_n686));
  NAND2_HPNW1  g0301(.A(new_n686), .B(new_n685), .Y(new_n687));
  NAND2_HPNW1  g0302(.A(\b[39] ), .B(\a[39] ), .Y(new_n688));
  NAND2_HPNW1  g0303(.A(new_n687), .B(new_n688), .Y(new_n689));
  XNOR2_HPNW1  g0304(.A(new_n684), .B(new_n689), .Y(\f[39] ));
  INV1_HPNW1   g0305(.A(new_n688), .Y(new_n691));
  AOI21_HPNW1  g0306(.A0(new_n687), .A1(new_n684), .B0(new_n691), .Y(new_n692));
  INV1_HPNW1   g0307(.A(\a[40] ), .Y(new_n693));
  INV1_HPNW1   g0308(.A(\b[40] ), .Y(new_n694));
  NAND2_HPNW1  g0309(.A(new_n694), .B(new_n693), .Y(new_n695));
  NAND2_HPNW1  g0310(.A(\b[40] ), .B(\a[40] ), .Y(new_n696));
  NAND2_HPNW1  g0311(.A(new_n695), .B(new_n696), .Y(new_n697));
  XOR2_HPNW1   g0312(.A(new_n697), .B(new_n692), .Y(\f[40] ));
  INV1_HPNW1   g0313(.A(new_n695), .Y(new_n699));
  OAI21_HPNW1  g0314(.A0(new_n699), .A1(new_n692), .B0(new_n696), .Y(new_n700));
  INV1_HPNW1   g0315(.A(\a[41] ), .Y(new_n701));
  INV1_HPNW1   g0316(.A(\b[41] ), .Y(new_n702));
  NAND2_HPNW1  g0317(.A(new_n702), .B(new_n701), .Y(new_n703));
  NAND2_HPNW1  g0318(.A(\b[41] ), .B(\a[41] ), .Y(new_n704));
  NAND2_HPNW1  g0319(.A(new_n703), .B(new_n704), .Y(new_n705));
  XNOR2_HPNW1  g0320(.A(new_n700), .B(new_n705), .Y(\f[41] ));
  INV1_HPNW1   g0321(.A(new_n704), .Y(new_n707));
  AOI21_HPNW1  g0322(.A0(new_n703), .A1(new_n700), .B0(new_n707), .Y(new_n708));
  INV1_HPNW1   g0323(.A(\a[42] ), .Y(new_n709));
  INV1_HPNW1   g0324(.A(\b[42] ), .Y(new_n710));
  NAND2_HPNW1  g0325(.A(new_n710), .B(new_n709), .Y(new_n711));
  NAND2_HPNW1  g0326(.A(\b[42] ), .B(\a[42] ), .Y(new_n712));
  NAND2_HPNW1  g0327(.A(new_n711), .B(new_n712), .Y(new_n713));
  XOR2_HPNW1   g0328(.A(new_n713), .B(new_n708), .Y(\f[42] ));
  INV1_HPNW1   g0329(.A(new_n711), .Y(new_n715));
  OAI21_HPNW1  g0330(.A0(new_n715), .A1(new_n708), .B0(new_n712), .Y(new_n716));
  INV1_HPNW1   g0331(.A(\a[43] ), .Y(new_n717));
  INV1_HPNW1   g0332(.A(\b[43] ), .Y(new_n718));
  NAND2_HPNW1  g0333(.A(new_n718), .B(new_n717), .Y(new_n719));
  NAND2_HPNW1  g0334(.A(\b[43] ), .B(\a[43] ), .Y(new_n720));
  NAND2_HPNW1  g0335(.A(new_n719), .B(new_n720), .Y(new_n721));
  XNOR2_HPNW1  g0336(.A(new_n716), .B(new_n721), .Y(\f[43] ));
  INV1_HPNW1   g0337(.A(new_n720), .Y(new_n723));
  AOI21_HPNW1  g0338(.A0(new_n719), .A1(new_n716), .B0(new_n723), .Y(new_n724));
  INV1_HPNW1   g0339(.A(\a[44] ), .Y(new_n725));
  INV1_HPNW1   g0340(.A(\b[44] ), .Y(new_n726));
  NAND2_HPNW1  g0341(.A(new_n726), .B(new_n725), .Y(new_n727));
  NAND2_HPNW1  g0342(.A(\b[44] ), .B(\a[44] ), .Y(new_n728));
  NAND2_HPNW1  g0343(.A(new_n727), .B(new_n728), .Y(new_n729));
  XOR2_HPNW1   g0344(.A(new_n729), .B(new_n724), .Y(\f[44] ));
  INV1_HPNW1   g0345(.A(new_n727), .Y(new_n731));
  OAI21_HPNW1  g0346(.A0(new_n731), .A1(new_n724), .B0(new_n728), .Y(new_n732));
  INV1_HPNW1   g0347(.A(\a[45] ), .Y(new_n733));
  INV1_HPNW1   g0348(.A(\b[45] ), .Y(new_n734));
  NAND2_HPNW1  g0349(.A(new_n734), .B(new_n733), .Y(new_n735));
  NAND2_HPNW1  g0350(.A(\b[45] ), .B(\a[45] ), .Y(new_n736));
  NAND2_HPNW1  g0351(.A(new_n735), .B(new_n736), .Y(new_n737));
  XNOR2_HPNW1  g0352(.A(new_n732), .B(new_n737), .Y(\f[45] ));
  INV1_HPNW1   g0353(.A(new_n736), .Y(new_n739));
  AOI21_HPNW1  g0354(.A0(new_n735), .A1(new_n732), .B0(new_n739), .Y(new_n740));
  INV1_HPNW1   g0355(.A(\a[46] ), .Y(new_n741));
  INV1_HPNW1   g0356(.A(\b[46] ), .Y(new_n742));
  NAND2_HPNW1  g0357(.A(new_n742), .B(new_n741), .Y(new_n743));
  NAND2_HPNW1  g0358(.A(\b[46] ), .B(\a[46] ), .Y(new_n744));
  NAND2_HPNW1  g0359(.A(new_n743), .B(new_n744), .Y(new_n745));
  XOR2_HPNW1   g0360(.A(new_n745), .B(new_n740), .Y(\f[46] ));
  INV1_HPNW1   g0361(.A(new_n743), .Y(new_n747));
  OAI21_HPNW1  g0362(.A0(new_n747), .A1(new_n740), .B0(new_n744), .Y(new_n748));
  INV1_HPNW1   g0363(.A(\a[47] ), .Y(new_n749));
  INV1_HPNW1   g0364(.A(\b[47] ), .Y(new_n750));
  NAND2_HPNW1  g0365(.A(new_n750), .B(new_n749), .Y(new_n751));
  NAND2_HPNW1  g0366(.A(\b[47] ), .B(\a[47] ), .Y(new_n752));
  NAND2_HPNW1  g0367(.A(new_n751), .B(new_n752), .Y(new_n753));
  XNOR2_HPNW1  g0368(.A(new_n748), .B(new_n753), .Y(\f[47] ));
  INV1_HPNW1   g0369(.A(new_n752), .Y(new_n755));
  AOI21_HPNW1  g0370(.A0(new_n751), .A1(new_n748), .B0(new_n755), .Y(new_n756));
  INV1_HPNW1   g0371(.A(\a[48] ), .Y(new_n757));
  INV1_HPNW1   g0372(.A(\b[48] ), .Y(new_n758));
  NAND2_HPNW1  g0373(.A(new_n758), .B(new_n757), .Y(new_n759));
  NAND2_HPNW1  g0374(.A(\b[48] ), .B(\a[48] ), .Y(new_n760));
  NAND2_HPNW1  g0375(.A(new_n759), .B(new_n760), .Y(new_n761));
  XOR2_HPNW1   g0376(.A(new_n761), .B(new_n756), .Y(\f[48] ));
  INV1_HPNW1   g0377(.A(new_n759), .Y(new_n763));
  OAI21_HPNW1  g0378(.A0(new_n763), .A1(new_n756), .B0(new_n760), .Y(new_n764));
  INV1_HPNW1   g0379(.A(\a[49] ), .Y(new_n765));
  INV1_HPNW1   g0380(.A(\b[49] ), .Y(new_n766));
  NAND2_HPNW1  g0381(.A(new_n766), .B(new_n765), .Y(new_n767));
  NAND2_HPNW1  g0382(.A(\b[49] ), .B(\a[49] ), .Y(new_n768));
  NAND2_HPNW1  g0383(.A(new_n767), .B(new_n768), .Y(new_n769));
  XNOR2_HPNW1  g0384(.A(new_n764), .B(new_n769), .Y(\f[49] ));
  INV1_HPNW1   g0385(.A(new_n768), .Y(new_n771));
  AOI21_HPNW1  g0386(.A0(new_n767), .A1(new_n764), .B0(new_n771), .Y(new_n772));
  INV1_HPNW1   g0387(.A(\a[50] ), .Y(new_n773));
  INV1_HPNW1   g0388(.A(\b[50] ), .Y(new_n774));
  NAND2_HPNW1  g0389(.A(new_n774), .B(new_n773), .Y(new_n775));
  NAND2_HPNW1  g0390(.A(\b[50] ), .B(\a[50] ), .Y(new_n776));
  NAND2_HPNW1  g0391(.A(new_n775), .B(new_n776), .Y(new_n777));
  XOR2_HPNW1   g0392(.A(new_n777), .B(new_n772), .Y(\f[50] ));
  INV1_HPNW1   g0393(.A(new_n775), .Y(new_n779));
  OAI21_HPNW1  g0394(.A0(new_n779), .A1(new_n772), .B0(new_n776), .Y(new_n780));
  INV1_HPNW1   g0395(.A(\a[51] ), .Y(new_n781));
  INV1_HPNW1   g0396(.A(\b[51] ), .Y(new_n782));
  NAND2_HPNW1  g0397(.A(new_n782), .B(new_n781), .Y(new_n783));
  NAND2_HPNW1  g0398(.A(\b[51] ), .B(\a[51] ), .Y(new_n784));
  NAND2_HPNW1  g0399(.A(new_n783), .B(new_n784), .Y(new_n785));
  XNOR2_HPNW1  g0400(.A(new_n780), .B(new_n785), .Y(\f[51] ));
  INV1_HPNW1   g0401(.A(new_n784), .Y(new_n787));
  AOI21_HPNW1  g0402(.A0(new_n783), .A1(new_n780), .B0(new_n787), .Y(new_n788));
  INV1_HPNW1   g0403(.A(\a[52] ), .Y(new_n789));
  INV1_HPNW1   g0404(.A(\b[52] ), .Y(new_n790));
  NAND2_HPNW1  g0405(.A(new_n790), .B(new_n789), .Y(new_n791));
  NAND2_HPNW1  g0406(.A(\b[52] ), .B(\a[52] ), .Y(new_n792));
  NAND2_HPNW1  g0407(.A(new_n791), .B(new_n792), .Y(new_n793));
  XOR2_HPNW1   g0408(.A(new_n793), .B(new_n788), .Y(\f[52] ));
  INV1_HPNW1   g0409(.A(new_n791), .Y(new_n795));
  OAI21_HPNW1  g0410(.A0(new_n795), .A1(new_n788), .B0(new_n792), .Y(new_n796));
  INV1_HPNW1   g0411(.A(\a[53] ), .Y(new_n797));
  INV1_HPNW1   g0412(.A(\b[53] ), .Y(new_n798));
  NAND2_HPNW1  g0413(.A(new_n798), .B(new_n797), .Y(new_n799));
  NAND2_HPNW1  g0414(.A(\b[53] ), .B(\a[53] ), .Y(new_n800));
  NAND2_HPNW1  g0415(.A(new_n799), .B(new_n800), .Y(new_n801));
  XNOR2_HPNW1  g0416(.A(new_n796), .B(new_n801), .Y(\f[53] ));
  INV1_HPNW1   g0417(.A(new_n800), .Y(new_n803));
  AOI21_HPNW1  g0418(.A0(new_n799), .A1(new_n796), .B0(new_n803), .Y(new_n804));
  INV1_HPNW1   g0419(.A(\a[54] ), .Y(new_n805));
  INV1_HPNW1   g0420(.A(\b[54] ), .Y(new_n806));
  NAND2_HPNW1  g0421(.A(new_n806), .B(new_n805), .Y(new_n807));
  NAND2_HPNW1  g0422(.A(\b[54] ), .B(\a[54] ), .Y(new_n808));
  NAND2_HPNW1  g0423(.A(new_n807), .B(new_n808), .Y(new_n809));
  XOR2_HPNW1   g0424(.A(new_n809), .B(new_n804), .Y(\f[54] ));
  INV1_HPNW1   g0425(.A(new_n807), .Y(new_n811));
  OAI21_HPNW1  g0426(.A0(new_n811), .A1(new_n804), .B0(new_n808), .Y(new_n812));
  INV1_HPNW1   g0427(.A(\a[55] ), .Y(new_n813));
  INV1_HPNW1   g0428(.A(\b[55] ), .Y(new_n814));
  NAND2_HPNW1  g0429(.A(new_n814), .B(new_n813), .Y(new_n815));
  NAND2_HPNW1  g0430(.A(\b[55] ), .B(\a[55] ), .Y(new_n816));
  NAND2_HPNW1  g0431(.A(new_n815), .B(new_n816), .Y(new_n817));
  XNOR2_HPNW1  g0432(.A(new_n812), .B(new_n817), .Y(\f[55] ));
  INV1_HPNW1   g0433(.A(new_n816), .Y(new_n819));
  AOI21_HPNW1  g0434(.A0(new_n815), .A1(new_n812), .B0(new_n819), .Y(new_n820));
  INV1_HPNW1   g0435(.A(\a[56] ), .Y(new_n821));
  INV1_HPNW1   g0436(.A(\b[56] ), .Y(new_n822));
  NAND2_HPNW1  g0437(.A(new_n822), .B(new_n821), .Y(new_n823));
  NAND2_HPNW1  g0438(.A(\b[56] ), .B(\a[56] ), .Y(new_n824));
  NAND2_HPNW1  g0439(.A(new_n823), .B(new_n824), .Y(new_n825));
  XOR2_HPNW1   g0440(.A(new_n825), .B(new_n820), .Y(\f[56] ));
  INV1_HPNW1   g0441(.A(new_n823), .Y(new_n827));
  OAI21_HPNW1  g0442(.A0(new_n827), .A1(new_n820), .B0(new_n824), .Y(new_n828));
  INV1_HPNW1   g0443(.A(\a[57] ), .Y(new_n829));
  INV1_HPNW1   g0444(.A(\b[57] ), .Y(new_n830));
  NAND2_HPNW1  g0445(.A(new_n830), .B(new_n829), .Y(new_n831));
  NAND2_HPNW1  g0446(.A(\b[57] ), .B(\a[57] ), .Y(new_n832));
  NAND2_HPNW1  g0447(.A(new_n831), .B(new_n832), .Y(new_n833));
  XNOR2_HPNW1  g0448(.A(new_n828), .B(new_n833), .Y(\f[57] ));
  INV1_HPNW1   g0449(.A(new_n832), .Y(new_n835));
  AOI21_HPNW1  g0450(.A0(new_n831), .A1(new_n828), .B0(new_n835), .Y(new_n836));
  INV1_HPNW1   g0451(.A(\a[58] ), .Y(new_n837));
  INV1_HPNW1   g0452(.A(\b[58] ), .Y(new_n838));
  NAND2_HPNW1  g0453(.A(new_n838), .B(new_n837), .Y(new_n839));
  NAND2_HPNW1  g0454(.A(\b[58] ), .B(\a[58] ), .Y(new_n840));
  NAND2_HPNW1  g0455(.A(new_n839), .B(new_n840), .Y(new_n841));
  XOR2_HPNW1   g0456(.A(new_n841), .B(new_n836), .Y(\f[58] ));
  INV1_HPNW1   g0457(.A(new_n839), .Y(new_n843));
  OAI21_HPNW1  g0458(.A0(new_n843), .A1(new_n836), .B0(new_n840), .Y(new_n844));
  INV1_HPNW1   g0459(.A(\a[59] ), .Y(new_n845));
  INV1_HPNW1   g0460(.A(\b[59] ), .Y(new_n846));
  NAND2_HPNW1  g0461(.A(new_n846), .B(new_n845), .Y(new_n847));
  NAND2_HPNW1  g0462(.A(\b[59] ), .B(\a[59] ), .Y(new_n848));
  NAND2_HPNW1  g0463(.A(new_n847), .B(new_n848), .Y(new_n849));
  XNOR2_HPNW1  g0464(.A(new_n844), .B(new_n849), .Y(\f[59] ));
  INV1_HPNW1   g0465(.A(new_n848), .Y(new_n851));
  AOI21_HPNW1  g0466(.A0(new_n847), .A1(new_n844), .B0(new_n851), .Y(new_n852));
  INV1_HPNW1   g0467(.A(\a[60] ), .Y(new_n853));
  INV1_HPNW1   g0468(.A(\b[60] ), .Y(new_n854));
  NAND2_HPNW1  g0469(.A(new_n854), .B(new_n853), .Y(new_n855));
  NAND2_HPNW1  g0470(.A(\b[60] ), .B(\a[60] ), .Y(new_n856));
  NAND2_HPNW1  g0471(.A(new_n855), .B(new_n856), .Y(new_n857));
  XOR2_HPNW1   g0472(.A(new_n857), .B(new_n852), .Y(\f[60] ));
  INV1_HPNW1   g0473(.A(new_n855), .Y(new_n859));
  OAI21_HPNW1  g0474(.A0(new_n859), .A1(new_n852), .B0(new_n856), .Y(new_n860));
  INV1_HPNW1   g0475(.A(\a[61] ), .Y(new_n861));
  INV1_HPNW1   g0476(.A(\b[61] ), .Y(new_n862));
  NAND2_HPNW1  g0477(.A(new_n862), .B(new_n861), .Y(new_n863));
  NAND2_HPNW1  g0478(.A(\b[61] ), .B(\a[61] ), .Y(new_n864));
  NAND2_HPNW1  g0479(.A(new_n863), .B(new_n864), .Y(new_n865));
  XNOR2_HPNW1  g0480(.A(new_n860), .B(new_n865), .Y(\f[61] ));
  INV1_HPNW1   g0481(.A(new_n864), .Y(new_n867));
  AOI21_HPNW1  g0482(.A0(new_n863), .A1(new_n860), .B0(new_n867), .Y(new_n868));
  INV1_HPNW1   g0483(.A(\a[62] ), .Y(new_n869));
  INV1_HPNW1   g0484(.A(\b[62] ), .Y(new_n870));
  NAND2_HPNW1  g0485(.A(new_n870), .B(new_n869), .Y(new_n871));
  NAND2_HPNW1  g0486(.A(\b[62] ), .B(\a[62] ), .Y(new_n872));
  NAND2_HPNW1  g0487(.A(new_n871), .B(new_n872), .Y(new_n873));
  XOR2_HPNW1   g0488(.A(new_n873), .B(new_n868), .Y(\f[62] ));
  INV1_HPNW1   g0489(.A(new_n871), .Y(new_n875));
  OAI21_HPNW1  g0490(.A0(new_n875), .A1(new_n868), .B0(new_n872), .Y(new_n876));
  INV1_HPNW1   g0491(.A(\a[63] ), .Y(new_n877));
  INV1_HPNW1   g0492(.A(\b[63] ), .Y(new_n878));
  NAND2_HPNW1  g0493(.A(new_n878), .B(new_n877), .Y(new_n879));
  NAND2_HPNW1  g0494(.A(\b[63] ), .B(\a[63] ), .Y(new_n880));
  NAND2_HPNW1  g0495(.A(new_n879), .B(new_n880), .Y(new_n881));
  XNOR2_HPNW1  g0496(.A(new_n876), .B(new_n881), .Y(\f[63] ));
  INV1_HPNW1   g0497(.A(new_n880), .Y(new_n883));
  AOI21_HPNW1  g0498(.A0(new_n879), .A1(new_n876), .B0(new_n883), .Y(new_n884));
  INV1_HPNW1   g0499(.A(\a[64] ), .Y(new_n885));
  INV1_HPNW1   g0500(.A(\b[64] ), .Y(new_n886));
  NAND2_HPNW1  g0501(.A(new_n886), .B(new_n885), .Y(new_n887));
  NAND2_HPNW1  g0502(.A(\b[64] ), .B(\a[64] ), .Y(new_n888));
  NAND2_HPNW1  g0503(.A(new_n887), .B(new_n888), .Y(new_n889));
  XOR2_HPNW1   g0504(.A(new_n889), .B(new_n884), .Y(\f[64] ));
  INV1_HPNW1   g0505(.A(new_n887), .Y(new_n891));
  OAI21_HPNW1  g0506(.A0(new_n891), .A1(new_n884), .B0(new_n888), .Y(new_n892));
  INV1_HPNW1   g0507(.A(\a[65] ), .Y(new_n893));
  INV1_HPNW1   g0508(.A(\b[65] ), .Y(new_n894));
  NAND2_HPNW1  g0509(.A(new_n894), .B(new_n893), .Y(new_n895));
  NAND2_HPNW1  g0510(.A(\b[65] ), .B(\a[65] ), .Y(new_n896));
  NAND2_HPNW1  g0511(.A(new_n895), .B(new_n896), .Y(new_n897));
  XNOR2_HPNW1  g0512(.A(new_n892), .B(new_n897), .Y(\f[65] ));
  INV1_HPNW1   g0513(.A(new_n896), .Y(new_n899));
  AOI21_HPNW1  g0514(.A0(new_n895), .A1(new_n892), .B0(new_n899), .Y(new_n900));
  INV1_HPNW1   g0515(.A(\a[66] ), .Y(new_n901));
  INV1_HPNW1   g0516(.A(\b[66] ), .Y(new_n902));
  NAND2_HPNW1  g0517(.A(new_n902), .B(new_n901), .Y(new_n903));
  NAND2_HPNW1  g0518(.A(\b[66] ), .B(\a[66] ), .Y(new_n904));
  NAND2_HPNW1  g0519(.A(new_n903), .B(new_n904), .Y(new_n905));
  XOR2_HPNW1   g0520(.A(new_n905), .B(new_n900), .Y(\f[66] ));
  INV1_HPNW1   g0521(.A(new_n903), .Y(new_n907));
  OAI21_HPNW1  g0522(.A0(new_n907), .A1(new_n900), .B0(new_n904), .Y(new_n908));
  INV1_HPNW1   g0523(.A(\a[67] ), .Y(new_n909));
  INV1_HPNW1   g0524(.A(\b[67] ), .Y(new_n910));
  NAND2_HPNW1  g0525(.A(new_n910), .B(new_n909), .Y(new_n911));
  NAND2_HPNW1  g0526(.A(\b[67] ), .B(\a[67] ), .Y(new_n912));
  NAND2_HPNW1  g0527(.A(new_n911), .B(new_n912), .Y(new_n913));
  XNOR2_HPNW1  g0528(.A(new_n908), .B(new_n913), .Y(\f[67] ));
  INV1_HPNW1   g0529(.A(new_n912), .Y(new_n915));
  AOI21_HPNW1  g0530(.A0(new_n911), .A1(new_n908), .B0(new_n915), .Y(new_n916));
  INV1_HPNW1   g0531(.A(\a[68] ), .Y(new_n917));
  INV1_HPNW1   g0532(.A(\b[68] ), .Y(new_n918));
  NAND2_HPNW1  g0533(.A(new_n918), .B(new_n917), .Y(new_n919));
  NAND2_HPNW1  g0534(.A(\b[68] ), .B(\a[68] ), .Y(new_n920));
  NAND2_HPNW1  g0535(.A(new_n919), .B(new_n920), .Y(new_n921));
  XOR2_HPNW1   g0536(.A(new_n921), .B(new_n916), .Y(\f[68] ));
  INV1_HPNW1   g0537(.A(new_n919), .Y(new_n923));
  OAI21_HPNW1  g0538(.A0(new_n923), .A1(new_n916), .B0(new_n920), .Y(new_n924));
  INV1_HPNW1   g0539(.A(\a[69] ), .Y(new_n925));
  INV1_HPNW1   g0540(.A(\b[69] ), .Y(new_n926));
  NAND2_HPNW1  g0541(.A(new_n926), .B(new_n925), .Y(new_n927));
  NAND2_HPNW1  g0542(.A(\b[69] ), .B(\a[69] ), .Y(new_n928));
  NAND2_HPNW1  g0543(.A(new_n927), .B(new_n928), .Y(new_n929));
  XNOR2_HPNW1  g0544(.A(new_n924), .B(new_n929), .Y(\f[69] ));
  INV1_HPNW1   g0545(.A(new_n928), .Y(new_n931));
  AOI21_HPNW1  g0546(.A0(new_n927), .A1(new_n924), .B0(new_n931), .Y(new_n932));
  INV1_HPNW1   g0547(.A(\a[70] ), .Y(new_n933));
  INV1_HPNW1   g0548(.A(\b[70] ), .Y(new_n934));
  NAND2_HPNW1  g0549(.A(new_n934), .B(new_n933), .Y(new_n935));
  NAND2_HPNW1  g0550(.A(\b[70] ), .B(\a[70] ), .Y(new_n936));
  NAND2_HPNW1  g0551(.A(new_n935), .B(new_n936), .Y(new_n937));
  XOR2_HPNW1   g0552(.A(new_n937), .B(new_n932), .Y(\f[70] ));
  INV1_HPNW1   g0553(.A(new_n935), .Y(new_n939));
  OAI21_HPNW1  g0554(.A0(new_n939), .A1(new_n932), .B0(new_n936), .Y(new_n940));
  INV1_HPNW1   g0555(.A(\a[71] ), .Y(new_n941));
  INV1_HPNW1   g0556(.A(\b[71] ), .Y(new_n942));
  NAND2_HPNW1  g0557(.A(new_n942), .B(new_n941), .Y(new_n943));
  NAND2_HPNW1  g0558(.A(\b[71] ), .B(\a[71] ), .Y(new_n944));
  NAND2_HPNW1  g0559(.A(new_n943), .B(new_n944), .Y(new_n945));
  XNOR2_HPNW1  g0560(.A(new_n940), .B(new_n945), .Y(\f[71] ));
  INV1_HPNW1   g0561(.A(new_n944), .Y(new_n947));
  AOI21_HPNW1  g0562(.A0(new_n943), .A1(new_n940), .B0(new_n947), .Y(new_n948));
  INV1_HPNW1   g0563(.A(\a[72] ), .Y(new_n949));
  INV1_HPNW1   g0564(.A(\b[72] ), .Y(new_n950));
  NAND2_HPNW1  g0565(.A(new_n950), .B(new_n949), .Y(new_n951));
  NAND2_HPNW1  g0566(.A(\b[72] ), .B(\a[72] ), .Y(new_n952));
  NAND2_HPNW1  g0567(.A(new_n951), .B(new_n952), .Y(new_n953));
  XOR2_HPNW1   g0568(.A(new_n953), .B(new_n948), .Y(\f[72] ));
  INV1_HPNW1   g0569(.A(new_n951), .Y(new_n955));
  OAI21_HPNW1  g0570(.A0(new_n955), .A1(new_n948), .B0(new_n952), .Y(new_n956));
  INV1_HPNW1   g0571(.A(\a[73] ), .Y(new_n957));
  INV1_HPNW1   g0572(.A(\b[73] ), .Y(new_n958));
  NAND2_HPNW1  g0573(.A(new_n958), .B(new_n957), .Y(new_n959));
  NAND2_HPNW1  g0574(.A(\b[73] ), .B(\a[73] ), .Y(new_n960));
  NAND2_HPNW1  g0575(.A(new_n959), .B(new_n960), .Y(new_n961));
  XNOR2_HPNW1  g0576(.A(new_n956), .B(new_n961), .Y(\f[73] ));
  INV1_HPNW1   g0577(.A(new_n960), .Y(new_n963));
  AOI21_HPNW1  g0578(.A0(new_n959), .A1(new_n956), .B0(new_n963), .Y(new_n964));
  INV1_HPNW1   g0579(.A(\a[74] ), .Y(new_n965));
  INV1_HPNW1   g0580(.A(\b[74] ), .Y(new_n966));
  NAND2_HPNW1  g0581(.A(new_n966), .B(new_n965), .Y(new_n967));
  NAND2_HPNW1  g0582(.A(\b[74] ), .B(\a[74] ), .Y(new_n968));
  NAND2_HPNW1  g0583(.A(new_n967), .B(new_n968), .Y(new_n969));
  XOR2_HPNW1   g0584(.A(new_n969), .B(new_n964), .Y(\f[74] ));
  INV1_HPNW1   g0585(.A(new_n967), .Y(new_n971));
  OAI21_HPNW1  g0586(.A0(new_n971), .A1(new_n964), .B0(new_n968), .Y(new_n972));
  INV1_HPNW1   g0587(.A(\a[75] ), .Y(new_n973));
  INV1_HPNW1   g0588(.A(\b[75] ), .Y(new_n974));
  NAND2_HPNW1  g0589(.A(new_n974), .B(new_n973), .Y(new_n975));
  NAND2_HPNW1  g0590(.A(\b[75] ), .B(\a[75] ), .Y(new_n976));
  NAND2_HPNW1  g0591(.A(new_n975), .B(new_n976), .Y(new_n977));
  XNOR2_HPNW1  g0592(.A(new_n972), .B(new_n977), .Y(\f[75] ));
  INV1_HPNW1   g0593(.A(new_n976), .Y(new_n979));
  AOI21_HPNW1  g0594(.A0(new_n975), .A1(new_n972), .B0(new_n979), .Y(new_n980));
  INV1_HPNW1   g0595(.A(\a[76] ), .Y(new_n981));
  INV1_HPNW1   g0596(.A(\b[76] ), .Y(new_n982));
  NAND2_HPNW1  g0597(.A(new_n982), .B(new_n981), .Y(new_n983));
  NAND2_HPNW1  g0598(.A(\b[76] ), .B(\a[76] ), .Y(new_n984));
  NAND2_HPNW1  g0599(.A(new_n983), .B(new_n984), .Y(new_n985));
  XOR2_HPNW1   g0600(.A(new_n985), .B(new_n980), .Y(\f[76] ));
  INV1_HPNW1   g0601(.A(new_n983), .Y(new_n987));
  OAI21_HPNW1  g0602(.A0(new_n987), .A1(new_n980), .B0(new_n984), .Y(new_n988));
  INV1_HPNW1   g0603(.A(\a[77] ), .Y(new_n989));
  INV1_HPNW1   g0604(.A(\b[77] ), .Y(new_n990));
  NAND2_HPNW1  g0605(.A(new_n990), .B(new_n989), .Y(new_n991));
  NAND2_HPNW1  g0606(.A(\b[77] ), .B(\a[77] ), .Y(new_n992));
  NAND2_HPNW1  g0607(.A(new_n991), .B(new_n992), .Y(new_n993));
  XNOR2_HPNW1  g0608(.A(new_n988), .B(new_n993), .Y(\f[77] ));
  INV1_HPNW1   g0609(.A(new_n992), .Y(new_n995));
  AOI21_HPNW1  g0610(.A0(new_n991), .A1(new_n988), .B0(new_n995), .Y(new_n996));
  INV1_HPNW1   g0611(.A(\a[78] ), .Y(new_n997));
  INV1_HPNW1   g0612(.A(\b[78] ), .Y(new_n998));
  NAND2_HPNW1  g0613(.A(new_n998), .B(new_n997), .Y(new_n999));
  NAND2_HPNW1  g0614(.A(\b[78] ), .B(\a[78] ), .Y(new_n1000));
  NAND2_HPNW1  g0615(.A(new_n999), .B(new_n1000), .Y(new_n1001));
  XOR2_HPNW1   g0616(.A(new_n1001), .B(new_n996), .Y(\f[78] ));
  INV1_HPNW1   g0617(.A(new_n999), .Y(new_n1003));
  OAI21_HPNW1  g0618(.A0(new_n1003), .A1(new_n996), .B0(new_n1000), .Y(new_n1004));
  INV1_HPNW1   g0619(.A(\a[79] ), .Y(new_n1005));
  INV1_HPNW1   g0620(.A(\b[79] ), .Y(new_n1006));
  NAND2_HPNW1  g0621(.A(new_n1006), .B(new_n1005), .Y(new_n1007));
  NAND2_HPNW1  g0622(.A(\b[79] ), .B(\a[79] ), .Y(new_n1008));
  NAND2_HPNW1  g0623(.A(new_n1007), .B(new_n1008), .Y(new_n1009));
  XNOR2_HPNW1  g0624(.A(new_n1004), .B(new_n1009), .Y(\f[79] ));
  INV1_HPNW1   g0625(.A(new_n1008), .Y(new_n1011));
  AOI21_HPNW1  g0626(.A0(new_n1007), .A1(new_n1004), .B0(new_n1011), .Y(new_n1012));
  INV1_HPNW1   g0627(.A(\a[80] ), .Y(new_n1013));
  INV1_HPNW1   g0628(.A(\b[80] ), .Y(new_n1014));
  NAND2_HPNW1  g0629(.A(new_n1014), .B(new_n1013), .Y(new_n1015));
  NAND2_HPNW1  g0630(.A(\b[80] ), .B(\a[80] ), .Y(new_n1016));
  NAND2_HPNW1  g0631(.A(new_n1015), .B(new_n1016), .Y(new_n1017));
  XOR2_HPNW1   g0632(.A(new_n1017), .B(new_n1012), .Y(\f[80] ));
  INV1_HPNW1   g0633(.A(new_n1015), .Y(new_n1019));
  OAI21_HPNW1  g0634(.A0(new_n1019), .A1(new_n1012), .B0(new_n1016), .Y(new_n1020));
  INV1_HPNW1   g0635(.A(\a[81] ), .Y(new_n1021));
  INV1_HPNW1   g0636(.A(\b[81] ), .Y(new_n1022));
  NAND2_HPNW1  g0637(.A(new_n1022), .B(new_n1021), .Y(new_n1023));
  NAND2_HPNW1  g0638(.A(\b[81] ), .B(\a[81] ), .Y(new_n1024));
  NAND2_HPNW1  g0639(.A(new_n1023), .B(new_n1024), .Y(new_n1025));
  XNOR2_HPNW1  g0640(.A(new_n1020), .B(new_n1025), .Y(\f[81] ));
  INV1_HPNW1   g0641(.A(new_n1024), .Y(new_n1027));
  AOI21_HPNW1  g0642(.A0(new_n1023), .A1(new_n1020), .B0(new_n1027), .Y(new_n1028));
  INV1_HPNW1   g0643(.A(\a[82] ), .Y(new_n1029));
  INV1_HPNW1   g0644(.A(\b[82] ), .Y(new_n1030));
  NAND2_HPNW1  g0645(.A(new_n1030), .B(new_n1029), .Y(new_n1031));
  NAND2_HPNW1  g0646(.A(\b[82] ), .B(\a[82] ), .Y(new_n1032));
  NAND2_HPNW1  g0647(.A(new_n1031), .B(new_n1032), .Y(new_n1033));
  XOR2_HPNW1   g0648(.A(new_n1033), .B(new_n1028), .Y(\f[82] ));
  INV1_HPNW1   g0649(.A(new_n1031), .Y(new_n1035));
  OAI21_HPNW1  g0650(.A0(new_n1035), .A1(new_n1028), .B0(new_n1032), .Y(new_n1036));
  INV1_HPNW1   g0651(.A(\a[83] ), .Y(new_n1037));
  INV1_HPNW1   g0652(.A(\b[83] ), .Y(new_n1038));
  NAND2_HPNW1  g0653(.A(new_n1038), .B(new_n1037), .Y(new_n1039));
  NAND2_HPNW1  g0654(.A(\b[83] ), .B(\a[83] ), .Y(new_n1040));
  NAND2_HPNW1  g0655(.A(new_n1039), .B(new_n1040), .Y(new_n1041));
  XNOR2_HPNW1  g0656(.A(new_n1036), .B(new_n1041), .Y(\f[83] ));
  INV1_HPNW1   g0657(.A(new_n1040), .Y(new_n1043));
  AOI21_HPNW1  g0658(.A0(new_n1039), .A1(new_n1036), .B0(new_n1043), .Y(new_n1044));
  INV1_HPNW1   g0659(.A(\a[84] ), .Y(new_n1045));
  INV1_HPNW1   g0660(.A(\b[84] ), .Y(new_n1046));
  NAND2_HPNW1  g0661(.A(new_n1046), .B(new_n1045), .Y(new_n1047));
  NAND2_HPNW1  g0662(.A(\b[84] ), .B(\a[84] ), .Y(new_n1048));
  NAND2_HPNW1  g0663(.A(new_n1047), .B(new_n1048), .Y(new_n1049));
  XOR2_HPNW1   g0664(.A(new_n1049), .B(new_n1044), .Y(\f[84] ));
  INV1_HPNW1   g0665(.A(new_n1047), .Y(new_n1051));
  OAI21_HPNW1  g0666(.A0(new_n1051), .A1(new_n1044), .B0(new_n1048), .Y(new_n1052));
  INV1_HPNW1   g0667(.A(\a[85] ), .Y(new_n1053));
  INV1_HPNW1   g0668(.A(\b[85] ), .Y(new_n1054));
  NAND2_HPNW1  g0669(.A(new_n1054), .B(new_n1053), .Y(new_n1055));
  NAND2_HPNW1  g0670(.A(\b[85] ), .B(\a[85] ), .Y(new_n1056));
  NAND2_HPNW1  g0671(.A(new_n1055), .B(new_n1056), .Y(new_n1057));
  XNOR2_HPNW1  g0672(.A(new_n1052), .B(new_n1057), .Y(\f[85] ));
  INV1_HPNW1   g0673(.A(new_n1056), .Y(new_n1059));
  AOI21_HPNW1  g0674(.A0(new_n1055), .A1(new_n1052), .B0(new_n1059), .Y(new_n1060));
  INV1_HPNW1   g0675(.A(\a[86] ), .Y(new_n1061));
  INV1_HPNW1   g0676(.A(\b[86] ), .Y(new_n1062));
  NAND2_HPNW1  g0677(.A(new_n1062), .B(new_n1061), .Y(new_n1063));
  NAND2_HPNW1  g0678(.A(\b[86] ), .B(\a[86] ), .Y(new_n1064));
  NAND2_HPNW1  g0679(.A(new_n1063), .B(new_n1064), .Y(new_n1065));
  XOR2_HPNW1   g0680(.A(new_n1065), .B(new_n1060), .Y(\f[86] ));
  INV1_HPNW1   g0681(.A(new_n1063), .Y(new_n1067));
  OAI21_HPNW1  g0682(.A0(new_n1067), .A1(new_n1060), .B0(new_n1064), .Y(new_n1068));
  INV1_HPNW1   g0683(.A(\a[87] ), .Y(new_n1069));
  INV1_HPNW1   g0684(.A(\b[87] ), .Y(new_n1070));
  NAND2_HPNW1  g0685(.A(new_n1070), .B(new_n1069), .Y(new_n1071));
  NAND2_HPNW1  g0686(.A(\b[87] ), .B(\a[87] ), .Y(new_n1072));
  NAND2_HPNW1  g0687(.A(new_n1071), .B(new_n1072), .Y(new_n1073));
  XNOR2_HPNW1  g0688(.A(new_n1068), .B(new_n1073), .Y(\f[87] ));
  INV1_HPNW1   g0689(.A(new_n1072), .Y(new_n1075));
  AOI21_HPNW1  g0690(.A0(new_n1071), .A1(new_n1068), .B0(new_n1075), .Y(new_n1076));
  INV1_HPNW1   g0691(.A(\a[88] ), .Y(new_n1077));
  INV1_HPNW1   g0692(.A(\b[88] ), .Y(new_n1078));
  NAND2_HPNW1  g0693(.A(new_n1078), .B(new_n1077), .Y(new_n1079));
  NAND2_HPNW1  g0694(.A(\b[88] ), .B(\a[88] ), .Y(new_n1080));
  NAND2_HPNW1  g0695(.A(new_n1079), .B(new_n1080), .Y(new_n1081));
  XOR2_HPNW1   g0696(.A(new_n1081), .B(new_n1076), .Y(\f[88] ));
  INV1_HPNW1   g0697(.A(new_n1079), .Y(new_n1083));
  OAI21_HPNW1  g0698(.A0(new_n1083), .A1(new_n1076), .B0(new_n1080), .Y(new_n1084));
  INV1_HPNW1   g0699(.A(\a[89] ), .Y(new_n1085));
  INV1_HPNW1   g0700(.A(\b[89] ), .Y(new_n1086));
  NAND2_HPNW1  g0701(.A(new_n1086), .B(new_n1085), .Y(new_n1087));
  NAND2_HPNW1  g0702(.A(\b[89] ), .B(\a[89] ), .Y(new_n1088));
  NAND2_HPNW1  g0703(.A(new_n1087), .B(new_n1088), .Y(new_n1089));
  XNOR2_HPNW1  g0704(.A(new_n1084), .B(new_n1089), .Y(\f[89] ));
  INV1_HPNW1   g0705(.A(new_n1088), .Y(new_n1091));
  AOI21_HPNW1  g0706(.A0(new_n1087), .A1(new_n1084), .B0(new_n1091), .Y(new_n1092));
  INV1_HPNW1   g0707(.A(\a[90] ), .Y(new_n1093));
  INV1_HPNW1   g0708(.A(\b[90] ), .Y(new_n1094));
  NAND2_HPNW1  g0709(.A(new_n1094), .B(new_n1093), .Y(new_n1095));
  NAND2_HPNW1  g0710(.A(\b[90] ), .B(\a[90] ), .Y(new_n1096));
  NAND2_HPNW1  g0711(.A(new_n1095), .B(new_n1096), .Y(new_n1097));
  XOR2_HPNW1   g0712(.A(new_n1097), .B(new_n1092), .Y(\f[90] ));
  INV1_HPNW1   g0713(.A(new_n1095), .Y(new_n1099));
  OAI21_HPNW1  g0714(.A0(new_n1099), .A1(new_n1092), .B0(new_n1096), .Y(new_n1100));
  INV1_HPNW1   g0715(.A(\a[91] ), .Y(new_n1101));
  INV1_HPNW1   g0716(.A(\b[91] ), .Y(new_n1102));
  NAND2_HPNW1  g0717(.A(new_n1102), .B(new_n1101), .Y(new_n1103));
  NAND2_HPNW1  g0718(.A(\b[91] ), .B(\a[91] ), .Y(new_n1104));
  NAND2_HPNW1  g0719(.A(new_n1103), .B(new_n1104), .Y(new_n1105));
  XNOR2_HPNW1  g0720(.A(new_n1100), .B(new_n1105), .Y(\f[91] ));
  INV1_HPNW1   g0721(.A(new_n1104), .Y(new_n1107));
  AOI21_HPNW1  g0722(.A0(new_n1103), .A1(new_n1100), .B0(new_n1107), .Y(new_n1108));
  INV1_HPNW1   g0723(.A(\a[92] ), .Y(new_n1109));
  INV1_HPNW1   g0724(.A(\b[92] ), .Y(new_n1110));
  NAND2_HPNW1  g0725(.A(new_n1110), .B(new_n1109), .Y(new_n1111));
  NAND2_HPNW1  g0726(.A(\b[92] ), .B(\a[92] ), .Y(new_n1112));
  NAND2_HPNW1  g0727(.A(new_n1111), .B(new_n1112), .Y(new_n1113));
  XOR2_HPNW1   g0728(.A(new_n1113), .B(new_n1108), .Y(\f[92] ));
  INV1_HPNW1   g0729(.A(new_n1111), .Y(new_n1115));
  OAI21_HPNW1  g0730(.A0(new_n1115), .A1(new_n1108), .B0(new_n1112), .Y(new_n1116));
  INV1_HPNW1   g0731(.A(\a[93] ), .Y(new_n1117));
  INV1_HPNW1   g0732(.A(\b[93] ), .Y(new_n1118));
  NAND2_HPNW1  g0733(.A(new_n1118), .B(new_n1117), .Y(new_n1119));
  NAND2_HPNW1  g0734(.A(\b[93] ), .B(\a[93] ), .Y(new_n1120));
  NAND2_HPNW1  g0735(.A(new_n1119), .B(new_n1120), .Y(new_n1121));
  XNOR2_HPNW1  g0736(.A(new_n1116), .B(new_n1121), .Y(\f[93] ));
  INV1_HPNW1   g0737(.A(new_n1120), .Y(new_n1123));
  AOI21_HPNW1  g0738(.A0(new_n1119), .A1(new_n1116), .B0(new_n1123), .Y(new_n1124));
  INV1_HPNW1   g0739(.A(\a[94] ), .Y(new_n1125));
  INV1_HPNW1   g0740(.A(\b[94] ), .Y(new_n1126));
  NAND2_HPNW1  g0741(.A(new_n1126), .B(new_n1125), .Y(new_n1127));
  NAND2_HPNW1  g0742(.A(\b[94] ), .B(\a[94] ), .Y(new_n1128));
  NAND2_HPNW1  g0743(.A(new_n1127), .B(new_n1128), .Y(new_n1129));
  XOR2_HPNW1   g0744(.A(new_n1129), .B(new_n1124), .Y(\f[94] ));
  INV1_HPNW1   g0745(.A(new_n1127), .Y(new_n1131));
  OAI21_HPNW1  g0746(.A0(new_n1131), .A1(new_n1124), .B0(new_n1128), .Y(new_n1132));
  INV1_HPNW1   g0747(.A(\a[95] ), .Y(new_n1133));
  INV1_HPNW1   g0748(.A(\b[95] ), .Y(new_n1134));
  NAND2_HPNW1  g0749(.A(new_n1134), .B(new_n1133), .Y(new_n1135));
  NAND2_HPNW1  g0750(.A(\b[95] ), .B(\a[95] ), .Y(new_n1136));
  NAND2_HPNW1  g0751(.A(new_n1135), .B(new_n1136), .Y(new_n1137));
  XNOR2_HPNW1  g0752(.A(new_n1132), .B(new_n1137), .Y(\f[95] ));
  INV1_HPNW1   g0753(.A(new_n1136), .Y(new_n1139));
  AOI21_HPNW1  g0754(.A0(new_n1135), .A1(new_n1132), .B0(new_n1139), .Y(new_n1140));
  INV1_HPNW1   g0755(.A(\a[96] ), .Y(new_n1141));
  INV1_HPNW1   g0756(.A(\b[96] ), .Y(new_n1142));
  NAND2_HPNW1  g0757(.A(new_n1142), .B(new_n1141), .Y(new_n1143));
  NAND2_HPNW1  g0758(.A(\b[96] ), .B(\a[96] ), .Y(new_n1144));
  NAND2_HPNW1  g0759(.A(new_n1143), .B(new_n1144), .Y(new_n1145));
  XOR2_HPNW1   g0760(.A(new_n1145), .B(new_n1140), .Y(\f[96] ));
  INV1_HPNW1   g0761(.A(new_n1143), .Y(new_n1147));
  OAI21_HPNW1  g0762(.A0(new_n1147), .A1(new_n1140), .B0(new_n1144), .Y(new_n1148));
  INV1_HPNW1   g0763(.A(\a[97] ), .Y(new_n1149));
  INV1_HPNW1   g0764(.A(\b[97] ), .Y(new_n1150));
  NAND2_HPNW1  g0765(.A(new_n1150), .B(new_n1149), .Y(new_n1151));
  NAND2_HPNW1  g0766(.A(\b[97] ), .B(\a[97] ), .Y(new_n1152));
  NAND2_HPNW1  g0767(.A(new_n1151), .B(new_n1152), .Y(new_n1153));
  XNOR2_HPNW1  g0768(.A(new_n1148), .B(new_n1153), .Y(\f[97] ));
  INV1_HPNW1   g0769(.A(new_n1152), .Y(new_n1155));
  AOI21_HPNW1  g0770(.A0(new_n1151), .A1(new_n1148), .B0(new_n1155), .Y(new_n1156));
  INV1_HPNW1   g0771(.A(\a[98] ), .Y(new_n1157));
  INV1_HPNW1   g0772(.A(\b[98] ), .Y(new_n1158));
  NAND2_HPNW1  g0773(.A(new_n1158), .B(new_n1157), .Y(new_n1159));
  NAND2_HPNW1  g0774(.A(\b[98] ), .B(\a[98] ), .Y(new_n1160));
  NAND2_HPNW1  g0775(.A(new_n1159), .B(new_n1160), .Y(new_n1161));
  XOR2_HPNW1   g0776(.A(new_n1161), .B(new_n1156), .Y(\f[98] ));
  INV1_HPNW1   g0777(.A(new_n1159), .Y(new_n1163));
  OAI21_HPNW1  g0778(.A0(new_n1163), .A1(new_n1156), .B0(new_n1160), .Y(new_n1164));
  INV1_HPNW1   g0779(.A(\a[99] ), .Y(new_n1165));
  INV1_HPNW1   g0780(.A(\b[99] ), .Y(new_n1166));
  NAND2_HPNW1  g0781(.A(new_n1166), .B(new_n1165), .Y(new_n1167));
  NAND2_HPNW1  g0782(.A(\b[99] ), .B(\a[99] ), .Y(new_n1168));
  NAND2_HPNW1  g0783(.A(new_n1167), .B(new_n1168), .Y(new_n1169));
  XNOR2_HPNW1  g0784(.A(new_n1164), .B(new_n1169), .Y(\f[99] ));
  INV1_HPNW1   g0785(.A(new_n1168), .Y(new_n1171));
  AOI21_HPNW1  g0786(.A0(new_n1167), .A1(new_n1164), .B0(new_n1171), .Y(new_n1172));
  INV1_HPNW1   g0787(.A(\a[100] ), .Y(new_n1173));
  INV1_HPNW1   g0788(.A(\b[100] ), .Y(new_n1174));
  NAND2_HPNW1  g0789(.A(new_n1174), .B(new_n1173), .Y(new_n1175));
  NAND2_HPNW1  g0790(.A(\b[100] ), .B(\a[100] ), .Y(new_n1176));
  NAND2_HPNW1  g0791(.A(new_n1175), .B(new_n1176), .Y(new_n1177));
  XOR2_HPNW1   g0792(.A(new_n1177), .B(new_n1172), .Y(\f[100] ));
  INV1_HPNW1   g0793(.A(new_n1175), .Y(new_n1179));
  OAI21_HPNW1  g0794(.A0(new_n1179), .A1(new_n1172), .B0(new_n1176), .Y(new_n1180));
  INV1_HPNW1   g0795(.A(\a[101] ), .Y(new_n1181));
  INV1_HPNW1   g0796(.A(\b[101] ), .Y(new_n1182));
  NAND2_HPNW1  g0797(.A(new_n1182), .B(new_n1181), .Y(new_n1183));
  NAND2_HPNW1  g0798(.A(\b[101] ), .B(\a[101] ), .Y(new_n1184));
  NAND2_HPNW1  g0799(.A(new_n1183), .B(new_n1184), .Y(new_n1185));
  XNOR2_HPNW1  g0800(.A(new_n1180), .B(new_n1185), .Y(\f[101] ));
  INV1_HPNW1   g0801(.A(new_n1184), .Y(new_n1187));
  AOI21_HPNW1  g0802(.A0(new_n1183), .A1(new_n1180), .B0(new_n1187), .Y(new_n1188));
  INV1_HPNW1   g0803(.A(\a[102] ), .Y(new_n1189));
  INV1_HPNW1   g0804(.A(\b[102] ), .Y(new_n1190));
  NAND2_HPNW1  g0805(.A(new_n1190), .B(new_n1189), .Y(new_n1191));
  NAND2_HPNW1  g0806(.A(\b[102] ), .B(\a[102] ), .Y(new_n1192));
  NAND2_HPNW1  g0807(.A(new_n1191), .B(new_n1192), .Y(new_n1193));
  XOR2_HPNW1   g0808(.A(new_n1193), .B(new_n1188), .Y(\f[102] ));
  INV1_HPNW1   g0809(.A(new_n1191), .Y(new_n1195));
  OAI21_HPNW1  g0810(.A0(new_n1195), .A1(new_n1188), .B0(new_n1192), .Y(new_n1196));
  INV1_HPNW1   g0811(.A(\a[103] ), .Y(new_n1197));
  INV1_HPNW1   g0812(.A(\b[103] ), .Y(new_n1198));
  NAND2_HPNW1  g0813(.A(new_n1198), .B(new_n1197), .Y(new_n1199));
  NAND2_HPNW1  g0814(.A(\b[103] ), .B(\a[103] ), .Y(new_n1200));
  NAND2_HPNW1  g0815(.A(new_n1199), .B(new_n1200), .Y(new_n1201));
  XNOR2_HPNW1  g0816(.A(new_n1196), .B(new_n1201), .Y(\f[103] ));
  INV1_HPNW1   g0817(.A(new_n1200), .Y(new_n1203));
  AOI21_HPNW1  g0818(.A0(new_n1199), .A1(new_n1196), .B0(new_n1203), .Y(new_n1204));
  INV1_HPNW1   g0819(.A(\a[104] ), .Y(new_n1205));
  INV1_HPNW1   g0820(.A(\b[104] ), .Y(new_n1206));
  NAND2_HPNW1  g0821(.A(new_n1206), .B(new_n1205), .Y(new_n1207));
  NAND2_HPNW1  g0822(.A(\b[104] ), .B(\a[104] ), .Y(new_n1208));
  NAND2_HPNW1  g0823(.A(new_n1207), .B(new_n1208), .Y(new_n1209));
  XOR2_HPNW1   g0824(.A(new_n1209), .B(new_n1204), .Y(\f[104] ));
  INV1_HPNW1   g0825(.A(new_n1207), .Y(new_n1211));
  OAI21_HPNW1  g0826(.A0(new_n1211), .A1(new_n1204), .B0(new_n1208), .Y(new_n1212));
  INV1_HPNW1   g0827(.A(\a[105] ), .Y(new_n1213));
  INV1_HPNW1   g0828(.A(\b[105] ), .Y(new_n1214));
  NAND2_HPNW1  g0829(.A(new_n1214), .B(new_n1213), .Y(new_n1215));
  NAND2_HPNW1  g0830(.A(\b[105] ), .B(\a[105] ), .Y(new_n1216));
  NAND2_HPNW1  g0831(.A(new_n1215), .B(new_n1216), .Y(new_n1217));
  XNOR2_HPNW1  g0832(.A(new_n1212), .B(new_n1217), .Y(\f[105] ));
  INV1_HPNW1   g0833(.A(new_n1216), .Y(new_n1219));
  AOI21_HPNW1  g0834(.A0(new_n1215), .A1(new_n1212), .B0(new_n1219), .Y(new_n1220));
  INV1_HPNW1   g0835(.A(\a[106] ), .Y(new_n1221));
  INV1_HPNW1   g0836(.A(\b[106] ), .Y(new_n1222));
  NAND2_HPNW1  g0837(.A(new_n1222), .B(new_n1221), .Y(new_n1223));
  NAND2_HPNW1  g0838(.A(\b[106] ), .B(\a[106] ), .Y(new_n1224));
  NAND2_HPNW1  g0839(.A(new_n1223), .B(new_n1224), .Y(new_n1225));
  XOR2_HPNW1   g0840(.A(new_n1225), .B(new_n1220), .Y(\f[106] ));
  INV1_HPNW1   g0841(.A(new_n1223), .Y(new_n1227));
  OAI21_HPNW1  g0842(.A0(new_n1227), .A1(new_n1220), .B0(new_n1224), .Y(new_n1228));
  INV1_HPNW1   g0843(.A(\a[107] ), .Y(new_n1229));
  INV1_HPNW1   g0844(.A(\b[107] ), .Y(new_n1230));
  NAND2_HPNW1  g0845(.A(new_n1230), .B(new_n1229), .Y(new_n1231));
  NAND2_HPNW1  g0846(.A(\b[107] ), .B(\a[107] ), .Y(new_n1232));
  NAND2_HPNW1  g0847(.A(new_n1231), .B(new_n1232), .Y(new_n1233));
  XNOR2_HPNW1  g0848(.A(new_n1228), .B(new_n1233), .Y(\f[107] ));
  INV1_HPNW1   g0849(.A(new_n1232), .Y(new_n1235));
  AOI21_HPNW1  g0850(.A0(new_n1231), .A1(new_n1228), .B0(new_n1235), .Y(new_n1236));
  INV1_HPNW1   g0851(.A(\a[108] ), .Y(new_n1237));
  INV1_HPNW1   g0852(.A(\b[108] ), .Y(new_n1238));
  NAND2_HPNW1  g0853(.A(new_n1238), .B(new_n1237), .Y(new_n1239));
  NAND2_HPNW1  g0854(.A(\b[108] ), .B(\a[108] ), .Y(new_n1240));
  NAND2_HPNW1  g0855(.A(new_n1239), .B(new_n1240), .Y(new_n1241));
  XOR2_HPNW1   g0856(.A(new_n1241), .B(new_n1236), .Y(\f[108] ));
  INV1_HPNW1   g0857(.A(new_n1239), .Y(new_n1243));
  OAI21_HPNW1  g0858(.A0(new_n1243), .A1(new_n1236), .B0(new_n1240), .Y(new_n1244));
  INV1_HPNW1   g0859(.A(\a[109] ), .Y(new_n1245));
  INV1_HPNW1   g0860(.A(\b[109] ), .Y(new_n1246));
  NAND2_HPNW1  g0861(.A(new_n1246), .B(new_n1245), .Y(new_n1247));
  NAND2_HPNW1  g0862(.A(\b[109] ), .B(\a[109] ), .Y(new_n1248));
  NAND2_HPNW1  g0863(.A(new_n1247), .B(new_n1248), .Y(new_n1249));
  XNOR2_HPNW1  g0864(.A(new_n1244), .B(new_n1249), .Y(\f[109] ));
  INV1_HPNW1   g0865(.A(new_n1248), .Y(new_n1251));
  AOI21_HPNW1  g0866(.A0(new_n1247), .A1(new_n1244), .B0(new_n1251), .Y(new_n1252));
  INV1_HPNW1   g0867(.A(\a[110] ), .Y(new_n1253));
  INV1_HPNW1   g0868(.A(\b[110] ), .Y(new_n1254));
  NAND2_HPNW1  g0869(.A(new_n1254), .B(new_n1253), .Y(new_n1255));
  NAND2_HPNW1  g0870(.A(\b[110] ), .B(\a[110] ), .Y(new_n1256));
  NAND2_HPNW1  g0871(.A(new_n1255), .B(new_n1256), .Y(new_n1257));
  XOR2_HPNW1   g0872(.A(new_n1257), .B(new_n1252), .Y(\f[110] ));
  INV1_HPNW1   g0873(.A(new_n1255), .Y(new_n1259));
  OAI21_HPNW1  g0874(.A0(new_n1259), .A1(new_n1252), .B0(new_n1256), .Y(new_n1260));
  INV1_HPNW1   g0875(.A(\a[111] ), .Y(new_n1261));
  INV1_HPNW1   g0876(.A(\b[111] ), .Y(new_n1262));
  NAND2_HPNW1  g0877(.A(new_n1262), .B(new_n1261), .Y(new_n1263));
  NAND2_HPNW1  g0878(.A(\b[111] ), .B(\a[111] ), .Y(new_n1264));
  NAND2_HPNW1  g0879(.A(new_n1263), .B(new_n1264), .Y(new_n1265));
  XNOR2_HPNW1  g0880(.A(new_n1260), .B(new_n1265), .Y(\f[111] ));
  INV1_HPNW1   g0881(.A(new_n1264), .Y(new_n1267));
  AOI21_HPNW1  g0882(.A0(new_n1263), .A1(new_n1260), .B0(new_n1267), .Y(new_n1268));
  INV1_HPNW1   g0883(.A(\a[112] ), .Y(new_n1269));
  INV1_HPNW1   g0884(.A(\b[112] ), .Y(new_n1270));
  NAND2_HPNW1  g0885(.A(new_n1270), .B(new_n1269), .Y(new_n1271));
  NAND2_HPNW1  g0886(.A(\b[112] ), .B(\a[112] ), .Y(new_n1272));
  NAND2_HPNW1  g0887(.A(new_n1271), .B(new_n1272), .Y(new_n1273));
  XOR2_HPNW1   g0888(.A(new_n1273), .B(new_n1268), .Y(\f[112] ));
  INV1_HPNW1   g0889(.A(new_n1271), .Y(new_n1275));
  OAI21_HPNW1  g0890(.A0(new_n1275), .A1(new_n1268), .B0(new_n1272), .Y(new_n1276));
  INV1_HPNW1   g0891(.A(\a[113] ), .Y(new_n1277));
  INV1_HPNW1   g0892(.A(\b[113] ), .Y(new_n1278));
  NAND2_HPNW1  g0893(.A(new_n1278), .B(new_n1277), .Y(new_n1279));
  NAND2_HPNW1  g0894(.A(\b[113] ), .B(\a[113] ), .Y(new_n1280));
  NAND2_HPNW1  g0895(.A(new_n1279), .B(new_n1280), .Y(new_n1281));
  XNOR2_HPNW1  g0896(.A(new_n1276), .B(new_n1281), .Y(\f[113] ));
  INV1_HPNW1   g0897(.A(new_n1280), .Y(new_n1283));
  AOI21_HPNW1  g0898(.A0(new_n1279), .A1(new_n1276), .B0(new_n1283), .Y(new_n1284));
  INV1_HPNW1   g0899(.A(\a[114] ), .Y(new_n1285));
  INV1_HPNW1   g0900(.A(\b[114] ), .Y(new_n1286));
  NAND2_HPNW1  g0901(.A(new_n1286), .B(new_n1285), .Y(new_n1287));
  NAND2_HPNW1  g0902(.A(\b[114] ), .B(\a[114] ), .Y(new_n1288));
  NAND2_HPNW1  g0903(.A(new_n1287), .B(new_n1288), .Y(new_n1289));
  XOR2_HPNW1   g0904(.A(new_n1289), .B(new_n1284), .Y(\f[114] ));
  INV1_HPNW1   g0905(.A(new_n1287), .Y(new_n1291));
  OAI21_HPNW1  g0906(.A0(new_n1291), .A1(new_n1284), .B0(new_n1288), .Y(new_n1292));
  INV1_HPNW1   g0907(.A(\a[115] ), .Y(new_n1293));
  INV1_HPNW1   g0908(.A(\b[115] ), .Y(new_n1294));
  NAND2_HPNW1  g0909(.A(new_n1294), .B(new_n1293), .Y(new_n1295));
  NAND2_HPNW1  g0910(.A(\b[115] ), .B(\a[115] ), .Y(new_n1296));
  NAND2_HPNW1  g0911(.A(new_n1295), .B(new_n1296), .Y(new_n1297));
  XNOR2_HPNW1  g0912(.A(new_n1292), .B(new_n1297), .Y(\f[115] ));
  INV1_HPNW1   g0913(.A(new_n1296), .Y(new_n1299));
  AOI21_HPNW1  g0914(.A0(new_n1295), .A1(new_n1292), .B0(new_n1299), .Y(new_n1300));
  INV1_HPNW1   g0915(.A(\a[116] ), .Y(new_n1301));
  INV1_HPNW1   g0916(.A(\b[116] ), .Y(new_n1302));
  NAND2_HPNW1  g0917(.A(new_n1302), .B(new_n1301), .Y(new_n1303));
  NAND2_HPNW1  g0918(.A(\b[116] ), .B(\a[116] ), .Y(new_n1304));
  NAND2_HPNW1  g0919(.A(new_n1303), .B(new_n1304), .Y(new_n1305));
  XOR2_HPNW1   g0920(.A(new_n1305), .B(new_n1300), .Y(\f[116] ));
  INV1_HPNW1   g0921(.A(new_n1303), .Y(new_n1307));
  OAI21_HPNW1  g0922(.A0(new_n1307), .A1(new_n1300), .B0(new_n1304), .Y(new_n1308));
  INV1_HPNW1   g0923(.A(\a[117] ), .Y(new_n1309));
  INV1_HPNW1   g0924(.A(\b[117] ), .Y(new_n1310));
  NAND2_HPNW1  g0925(.A(new_n1310), .B(new_n1309), .Y(new_n1311));
  NAND2_HPNW1  g0926(.A(\b[117] ), .B(\a[117] ), .Y(new_n1312));
  NAND2_HPNW1  g0927(.A(new_n1311), .B(new_n1312), .Y(new_n1313));
  XNOR2_HPNW1  g0928(.A(new_n1308), .B(new_n1313), .Y(\f[117] ));
  INV1_HPNW1   g0929(.A(new_n1312), .Y(new_n1315));
  AOI21_HPNW1  g0930(.A0(new_n1311), .A1(new_n1308), .B0(new_n1315), .Y(new_n1316));
  INV1_HPNW1   g0931(.A(\a[118] ), .Y(new_n1317));
  INV1_HPNW1   g0932(.A(\b[118] ), .Y(new_n1318));
  NAND2_HPNW1  g0933(.A(new_n1318), .B(new_n1317), .Y(new_n1319));
  NAND2_HPNW1  g0934(.A(\b[118] ), .B(\a[118] ), .Y(new_n1320));
  NAND2_HPNW1  g0935(.A(new_n1319), .B(new_n1320), .Y(new_n1321));
  XOR2_HPNW1   g0936(.A(new_n1321), .B(new_n1316), .Y(\f[118] ));
  INV1_HPNW1   g0937(.A(new_n1319), .Y(new_n1323));
  OAI21_HPNW1  g0938(.A0(new_n1323), .A1(new_n1316), .B0(new_n1320), .Y(new_n1324));
  INV1_HPNW1   g0939(.A(\a[119] ), .Y(new_n1325));
  INV1_HPNW1   g0940(.A(\b[119] ), .Y(new_n1326));
  NAND2_HPNW1  g0941(.A(new_n1326), .B(new_n1325), .Y(new_n1327));
  NAND2_HPNW1  g0942(.A(\b[119] ), .B(\a[119] ), .Y(new_n1328));
  NAND2_HPNW1  g0943(.A(new_n1327), .B(new_n1328), .Y(new_n1329));
  XNOR2_HPNW1  g0944(.A(new_n1324), .B(new_n1329), .Y(\f[119] ));
  INV1_HPNW1   g0945(.A(new_n1328), .Y(new_n1331));
  AOI21_HPNW1  g0946(.A0(new_n1327), .A1(new_n1324), .B0(new_n1331), .Y(new_n1332));
  INV1_HPNW1   g0947(.A(\a[120] ), .Y(new_n1333));
  INV1_HPNW1   g0948(.A(\b[120] ), .Y(new_n1334));
  NAND2_HPNW1  g0949(.A(new_n1334), .B(new_n1333), .Y(new_n1335));
  NAND2_HPNW1  g0950(.A(\b[120] ), .B(\a[120] ), .Y(new_n1336));
  NAND2_HPNW1  g0951(.A(new_n1335), .B(new_n1336), .Y(new_n1337));
  XOR2_HPNW1   g0952(.A(new_n1337), .B(new_n1332), .Y(\f[120] ));
  INV1_HPNW1   g0953(.A(new_n1335), .Y(new_n1339));
  OAI21_HPNW1  g0954(.A0(new_n1339), .A1(new_n1332), .B0(new_n1336), .Y(new_n1340));
  INV1_HPNW1   g0955(.A(\a[121] ), .Y(new_n1341));
  INV1_HPNW1   g0956(.A(\b[121] ), .Y(new_n1342));
  NAND2_HPNW1  g0957(.A(new_n1342), .B(new_n1341), .Y(new_n1343));
  NAND2_HPNW1  g0958(.A(\b[121] ), .B(\a[121] ), .Y(new_n1344));
  NAND2_HPNW1  g0959(.A(new_n1343), .B(new_n1344), .Y(new_n1345));
  XNOR2_HPNW1  g0960(.A(new_n1340), .B(new_n1345), .Y(\f[121] ));
  INV1_HPNW1   g0961(.A(new_n1344), .Y(new_n1347));
  AOI21_HPNW1  g0962(.A0(new_n1343), .A1(new_n1340), .B0(new_n1347), .Y(new_n1348));
  INV1_HPNW1   g0963(.A(\a[122] ), .Y(new_n1349));
  INV1_HPNW1   g0964(.A(\b[122] ), .Y(new_n1350));
  NAND2_HPNW1  g0965(.A(new_n1350), .B(new_n1349), .Y(new_n1351));
  NAND2_HPNW1  g0966(.A(\b[122] ), .B(\a[122] ), .Y(new_n1352));
  NAND2_HPNW1  g0967(.A(new_n1351), .B(new_n1352), .Y(new_n1353));
  XOR2_HPNW1   g0968(.A(new_n1353), .B(new_n1348), .Y(\f[122] ));
  INV1_HPNW1   g0969(.A(new_n1351), .Y(new_n1355));
  OAI21_HPNW1  g0970(.A0(new_n1355), .A1(new_n1348), .B0(new_n1352), .Y(new_n1356));
  INV1_HPNW1   g0971(.A(\a[123] ), .Y(new_n1357));
  INV1_HPNW1   g0972(.A(\b[123] ), .Y(new_n1358));
  NAND2_HPNW1  g0973(.A(new_n1358), .B(new_n1357), .Y(new_n1359));
  NAND2_HPNW1  g0974(.A(\b[123] ), .B(\a[123] ), .Y(new_n1360));
  NAND2_HPNW1  g0975(.A(new_n1359), .B(new_n1360), .Y(new_n1361));
  XNOR2_HPNW1  g0976(.A(new_n1356), .B(new_n1361), .Y(\f[123] ));
  INV1_HPNW1   g0977(.A(new_n1360), .Y(new_n1363));
  AOI21_HPNW1  g0978(.A0(new_n1359), .A1(new_n1356), .B0(new_n1363), .Y(new_n1364));
  INV1_HPNW1   g0979(.A(\a[124] ), .Y(new_n1365));
  INV1_HPNW1   g0980(.A(\b[124] ), .Y(new_n1366));
  NAND2_HPNW1  g0981(.A(new_n1366), .B(new_n1365), .Y(new_n1367));
  NAND2_HPNW1  g0982(.A(\b[124] ), .B(\a[124] ), .Y(new_n1368));
  NAND2_HPNW1  g0983(.A(new_n1367), .B(new_n1368), .Y(new_n1369));
  XOR2_HPNW1   g0984(.A(new_n1369), .B(new_n1364), .Y(\f[124] ));
  INV1_HPNW1   g0985(.A(new_n1367), .Y(new_n1371));
  OAI21_HPNW1  g0986(.A0(new_n1371), .A1(new_n1364), .B0(new_n1368), .Y(new_n1372));
  INV1_HPNW1   g0987(.A(\a[125] ), .Y(new_n1373));
  INV1_HPNW1   g0988(.A(\b[125] ), .Y(new_n1374));
  NAND2_HPNW1  g0989(.A(new_n1374), .B(new_n1373), .Y(new_n1375));
  NAND2_HPNW1  g0990(.A(\b[125] ), .B(\a[125] ), .Y(new_n1376));
  NAND2_HPNW1  g0991(.A(new_n1375), .B(new_n1376), .Y(new_n1377));
  XNOR2_HPNW1  g0992(.A(new_n1372), .B(new_n1377), .Y(\f[125] ));
  NAND2_HPNW1  g0993(.A(new_n1372), .B(new_n1375), .Y(new_n1379));
  NAND2_HPNW1  g0994(.A(new_n1379), .B(new_n1376), .Y(new_n1380));
  INV1_HPNW1   g0995(.A(\a[126] ), .Y(new_n1381));
  INV1_HPNW1   g0996(.A(\b[126] ), .Y(new_n1382));
  NAND2_HPNW1  g0997(.A(new_n1382), .B(new_n1381), .Y(new_n1383));
  NAND2_HPNW1  g0998(.A(\b[126] ), .B(\a[126] ), .Y(new_n1384));
  AOI21_HPNW1  g0999(.A0(new_n1384), .A1(new_n1383), .B0(new_n1380), .Y(new_n1385));
  INV1_HPNW1   g1000(.A(new_n1376), .Y(new_n1386));
  AOI21_HPNW1  g1001(.A0(new_n1375), .A1(new_n1372), .B0(new_n1386), .Y(new_n1387));
  NAND2_HPNW1  g1002(.A(new_n1383), .B(new_n1384), .Y(new_n1388));
  NOR2_HPNW1   g1003(.A(new_n1388), .B(new_n1387), .Y(new_n1389));
  NOR2_HPNW1   g1004(.A(new_n1389), .B(new_n1385), .Y(\f[126] ));
  INV1_HPNW1   g1005(.A(new_n1383), .Y(new_n1391));
  OAI21_HPNW1  g1006(.A0(new_n1391), .A1(new_n1387), .B0(new_n1384), .Y(new_n1392));
  XOR2_HPNW1   g1007(.A(\b[127] ), .B(\a[127] ), .Y(new_n1393));
  NOR2_HPNW1   g1008(.A(new_n1393), .B(new_n1392), .Y(new_n1394));
  OAI21_HPNW1  g1009(.A0(new_n390), .A1(new_n392), .B0(new_n394), .Y(new_n1395));
  INV1_HPNW1   g1010(.A(new_n402), .Y(new_n1396));
  AOI21_HPNW1  g1011(.A0(new_n395), .A1(new_n1395), .B0(new_n1396), .Y(new_n1397));
  OAI21_HPNW1  g1012(.A0(new_n406), .A1(new_n1397), .B0(new_n409), .Y(new_n1398));
  AOI21_HPNW1  g1013(.A0(new_n410), .A1(new_n1398), .B0(new_n414), .Y(new_n1399));
  OAI21_HPNW1  g1014(.A0(new_n419), .A1(new_n1399), .B0(new_n423), .Y(new_n1400));
  INV1_HPNW1   g1015(.A(new_n431), .Y(new_n1401));
  AOI21_HPNW1  g1016(.A0(new_n424), .A1(new_n1400), .B0(new_n1401), .Y(new_n1402));
  OAI21_HPNW1  g1017(.A0(new_n435), .A1(new_n1402), .B0(new_n439), .Y(new_n1403));
  INV1_HPNW1   g1018(.A(new_n447), .Y(new_n1404));
  AOI21_HPNW1  g1019(.A0(new_n440), .A1(new_n1403), .B0(new_n1404), .Y(new_n1405));
  OAI21_HPNW1  g1020(.A0(new_n451), .A1(new_n1405), .B0(new_n455), .Y(new_n1406));
  INV1_HPNW1   g1021(.A(new_n463), .Y(new_n1407));
  AOI21_HPNW1  g1022(.A0(new_n456), .A1(new_n1406), .B0(new_n1407), .Y(new_n1408));
  OAI21_HPNW1  g1023(.A0(new_n467), .A1(new_n1408), .B0(new_n471), .Y(new_n1409));
  INV1_HPNW1   g1024(.A(new_n479), .Y(new_n1410));
  AOI21_HPNW1  g1025(.A0(new_n472), .A1(new_n1409), .B0(new_n1410), .Y(new_n1411));
  OAI21_HPNW1  g1026(.A0(new_n483), .A1(new_n1411), .B0(new_n487), .Y(new_n1412));
  INV1_HPNW1   g1027(.A(new_n495), .Y(new_n1413));
  AOI21_HPNW1  g1028(.A0(new_n488), .A1(new_n1412), .B0(new_n1413), .Y(new_n1414));
  OAI21_HPNW1  g1029(.A0(new_n499), .A1(new_n1414), .B0(new_n503), .Y(new_n1415));
  INV1_HPNW1   g1030(.A(new_n511), .Y(new_n1416));
  AOI21_HPNW1  g1031(.A0(new_n504), .A1(new_n1415), .B0(new_n1416), .Y(new_n1417));
  OAI21_HPNW1  g1032(.A0(new_n515), .A1(new_n1417), .B0(new_n519), .Y(new_n1418));
  INV1_HPNW1   g1033(.A(new_n527), .Y(new_n1419));
  AOI21_HPNW1  g1034(.A0(new_n520), .A1(new_n1418), .B0(new_n1419), .Y(new_n1420));
  OAI21_HPNW1  g1035(.A0(new_n531), .A1(new_n1420), .B0(new_n535), .Y(new_n1421));
  INV1_HPNW1   g1036(.A(new_n543), .Y(new_n1422));
  AOI21_HPNW1  g1037(.A0(new_n536), .A1(new_n1421), .B0(new_n1422), .Y(new_n1423));
  OAI21_HPNW1  g1038(.A0(new_n547), .A1(new_n1423), .B0(new_n551), .Y(new_n1424));
  INV1_HPNW1   g1039(.A(new_n559), .Y(new_n1425));
  AOI21_HPNW1  g1040(.A0(new_n552), .A1(new_n1424), .B0(new_n1425), .Y(new_n1426));
  OAI21_HPNW1  g1041(.A0(new_n563), .A1(new_n1426), .B0(new_n567), .Y(new_n1427));
  INV1_HPNW1   g1042(.A(new_n575), .Y(new_n1428));
  AOI21_HPNW1  g1043(.A0(new_n568), .A1(new_n1427), .B0(new_n1428), .Y(new_n1429));
  OAI21_HPNW1  g1044(.A0(new_n579), .A1(new_n1429), .B0(new_n583), .Y(new_n1430));
  INV1_HPNW1   g1045(.A(new_n591), .Y(new_n1431));
  AOI21_HPNW1  g1046(.A0(new_n584), .A1(new_n1430), .B0(new_n1431), .Y(new_n1432));
  OAI21_HPNW1  g1047(.A0(new_n595), .A1(new_n1432), .B0(new_n599), .Y(new_n1433));
  INV1_HPNW1   g1048(.A(new_n607), .Y(new_n1434));
  AOI21_HPNW1  g1049(.A0(new_n600), .A1(new_n1433), .B0(new_n1434), .Y(new_n1435));
  OAI21_HPNW1  g1050(.A0(new_n611), .A1(new_n1435), .B0(new_n615), .Y(new_n1436));
  INV1_HPNW1   g1051(.A(new_n623), .Y(new_n1437));
  AOI21_HPNW1  g1052(.A0(new_n616), .A1(new_n1436), .B0(new_n1437), .Y(new_n1438));
  OAI21_HPNW1  g1053(.A0(new_n627), .A1(new_n1438), .B0(new_n631), .Y(new_n1439));
  INV1_HPNW1   g1054(.A(new_n639), .Y(new_n1440));
  AOI21_HPNW1  g1055(.A0(new_n632), .A1(new_n1439), .B0(new_n1440), .Y(new_n1441));
  OAI21_HPNW1  g1056(.A0(new_n643), .A1(new_n1441), .B0(new_n647), .Y(new_n1442));
  INV1_HPNW1   g1057(.A(new_n655), .Y(new_n1443));
  AOI21_HPNW1  g1058(.A0(new_n648), .A1(new_n1442), .B0(new_n1443), .Y(new_n1444));
  OAI21_HPNW1  g1059(.A0(new_n659), .A1(new_n1444), .B0(new_n663), .Y(new_n1445));
  INV1_HPNW1   g1060(.A(new_n671), .Y(new_n1446));
  AOI21_HPNW1  g1061(.A0(new_n664), .A1(new_n1445), .B0(new_n1446), .Y(new_n1447));
  OAI21_HPNW1  g1062(.A0(new_n675), .A1(new_n1447), .B0(new_n679), .Y(new_n1448));
  INV1_HPNW1   g1063(.A(new_n687), .Y(new_n1449));
  AOI21_HPNW1  g1064(.A0(new_n680), .A1(new_n1448), .B0(new_n1449), .Y(new_n1450));
  OAI21_HPNW1  g1065(.A0(new_n691), .A1(new_n1450), .B0(new_n695), .Y(new_n1451));
  INV1_HPNW1   g1066(.A(new_n703), .Y(new_n1452));
  AOI21_HPNW1  g1067(.A0(new_n696), .A1(new_n1451), .B0(new_n1452), .Y(new_n1453));
  OAI21_HPNW1  g1068(.A0(new_n707), .A1(new_n1453), .B0(new_n711), .Y(new_n1454));
  INV1_HPNW1   g1069(.A(new_n719), .Y(new_n1455));
  AOI21_HPNW1  g1070(.A0(new_n712), .A1(new_n1454), .B0(new_n1455), .Y(new_n1456));
  OAI21_HPNW1  g1071(.A0(new_n723), .A1(new_n1456), .B0(new_n727), .Y(new_n1457));
  INV1_HPNW1   g1072(.A(new_n735), .Y(new_n1458));
  AOI21_HPNW1  g1073(.A0(new_n728), .A1(new_n1457), .B0(new_n1458), .Y(new_n1459));
  OAI21_HPNW1  g1074(.A0(new_n739), .A1(new_n1459), .B0(new_n743), .Y(new_n1460));
  INV1_HPNW1   g1075(.A(new_n751), .Y(new_n1461));
  AOI21_HPNW1  g1076(.A0(new_n744), .A1(new_n1460), .B0(new_n1461), .Y(new_n1462));
  OAI21_HPNW1  g1077(.A0(new_n755), .A1(new_n1462), .B0(new_n759), .Y(new_n1463));
  INV1_HPNW1   g1078(.A(new_n767), .Y(new_n1464));
  AOI21_HPNW1  g1079(.A0(new_n760), .A1(new_n1463), .B0(new_n1464), .Y(new_n1465));
  OAI21_HPNW1  g1080(.A0(new_n771), .A1(new_n1465), .B0(new_n775), .Y(new_n1466));
  INV1_HPNW1   g1081(.A(new_n783), .Y(new_n1467));
  AOI21_HPNW1  g1082(.A0(new_n776), .A1(new_n1466), .B0(new_n1467), .Y(new_n1468));
  OAI21_HPNW1  g1083(.A0(new_n787), .A1(new_n1468), .B0(new_n791), .Y(new_n1469));
  INV1_HPNW1   g1084(.A(new_n799), .Y(new_n1470));
  AOI21_HPNW1  g1085(.A0(new_n792), .A1(new_n1469), .B0(new_n1470), .Y(new_n1471));
  OAI21_HPNW1  g1086(.A0(new_n803), .A1(new_n1471), .B0(new_n807), .Y(new_n1472));
  INV1_HPNW1   g1087(.A(new_n815), .Y(new_n1473));
  AOI21_HPNW1  g1088(.A0(new_n808), .A1(new_n1472), .B0(new_n1473), .Y(new_n1474));
  OAI21_HPNW1  g1089(.A0(new_n819), .A1(new_n1474), .B0(new_n823), .Y(new_n1475));
  INV1_HPNW1   g1090(.A(new_n831), .Y(new_n1476));
  AOI21_HPNW1  g1091(.A0(new_n824), .A1(new_n1475), .B0(new_n1476), .Y(new_n1477));
  OAI21_HPNW1  g1092(.A0(new_n835), .A1(new_n1477), .B0(new_n839), .Y(new_n1478));
  INV1_HPNW1   g1093(.A(new_n847), .Y(new_n1479));
  AOI21_HPNW1  g1094(.A0(new_n840), .A1(new_n1478), .B0(new_n1479), .Y(new_n1480));
  OAI21_HPNW1  g1095(.A0(new_n851), .A1(new_n1480), .B0(new_n855), .Y(new_n1481));
  INV1_HPNW1   g1096(.A(new_n863), .Y(new_n1482));
  AOI21_HPNW1  g1097(.A0(new_n856), .A1(new_n1481), .B0(new_n1482), .Y(new_n1483));
  OAI21_HPNW1  g1098(.A0(new_n867), .A1(new_n1483), .B0(new_n871), .Y(new_n1484));
  INV1_HPNW1   g1099(.A(new_n879), .Y(new_n1485));
  AOI21_HPNW1  g1100(.A0(new_n872), .A1(new_n1484), .B0(new_n1485), .Y(new_n1486));
  OAI21_HPNW1  g1101(.A0(new_n883), .A1(new_n1486), .B0(new_n887), .Y(new_n1487));
  INV1_HPNW1   g1102(.A(new_n895), .Y(new_n1488));
  AOI21_HPNW1  g1103(.A0(new_n888), .A1(new_n1487), .B0(new_n1488), .Y(new_n1489));
  OAI21_HPNW1  g1104(.A0(new_n899), .A1(new_n1489), .B0(new_n903), .Y(new_n1490));
  INV1_HPNW1   g1105(.A(new_n911), .Y(new_n1491));
  AOI21_HPNW1  g1106(.A0(new_n904), .A1(new_n1490), .B0(new_n1491), .Y(new_n1492));
  OAI21_HPNW1  g1107(.A0(new_n915), .A1(new_n1492), .B0(new_n919), .Y(new_n1493));
  INV1_HPNW1   g1108(.A(new_n927), .Y(new_n1494));
  AOI21_HPNW1  g1109(.A0(new_n920), .A1(new_n1493), .B0(new_n1494), .Y(new_n1495));
  OAI21_HPNW1  g1110(.A0(new_n931), .A1(new_n1495), .B0(new_n935), .Y(new_n1496));
  INV1_HPNW1   g1111(.A(new_n943), .Y(new_n1497));
  AOI21_HPNW1  g1112(.A0(new_n936), .A1(new_n1496), .B0(new_n1497), .Y(new_n1498));
  OAI21_HPNW1  g1113(.A0(new_n947), .A1(new_n1498), .B0(new_n951), .Y(new_n1499));
  INV1_HPNW1   g1114(.A(new_n959), .Y(new_n1500));
  AOI21_HPNW1  g1115(.A0(new_n952), .A1(new_n1499), .B0(new_n1500), .Y(new_n1501));
  OAI21_HPNW1  g1116(.A0(new_n963), .A1(new_n1501), .B0(new_n967), .Y(new_n1502));
  INV1_HPNW1   g1117(.A(new_n975), .Y(new_n1503));
  AOI21_HPNW1  g1118(.A0(new_n968), .A1(new_n1502), .B0(new_n1503), .Y(new_n1504));
  OAI21_HPNW1  g1119(.A0(new_n979), .A1(new_n1504), .B0(new_n983), .Y(new_n1505));
  INV1_HPNW1   g1120(.A(new_n991), .Y(new_n1506));
  AOI21_HPNW1  g1121(.A0(new_n984), .A1(new_n1505), .B0(new_n1506), .Y(new_n1507));
  OAI21_HPNW1  g1122(.A0(new_n995), .A1(new_n1507), .B0(new_n999), .Y(new_n1508));
  INV1_HPNW1   g1123(.A(new_n1007), .Y(new_n1509));
  AOI21_HPNW1  g1124(.A0(new_n1000), .A1(new_n1508), .B0(new_n1509), .Y(new_n1510));
  OAI21_HPNW1  g1125(.A0(new_n1011), .A1(new_n1510), .B0(new_n1015), .Y(new_n1511));
  INV1_HPNW1   g1126(.A(new_n1023), .Y(new_n1512));
  AOI21_HPNW1  g1127(.A0(new_n1016), .A1(new_n1511), .B0(new_n1512), .Y(new_n1513));
  OAI21_HPNW1  g1128(.A0(new_n1027), .A1(new_n1513), .B0(new_n1031), .Y(new_n1514));
  INV1_HPNW1   g1129(.A(new_n1039), .Y(new_n1515));
  AOI21_HPNW1  g1130(.A0(new_n1032), .A1(new_n1514), .B0(new_n1515), .Y(new_n1516));
  OAI21_HPNW1  g1131(.A0(new_n1043), .A1(new_n1516), .B0(new_n1047), .Y(new_n1517));
  INV1_HPNW1   g1132(.A(new_n1055), .Y(new_n1518));
  AOI21_HPNW1  g1133(.A0(new_n1048), .A1(new_n1517), .B0(new_n1518), .Y(new_n1519));
  OAI21_HPNW1  g1134(.A0(new_n1059), .A1(new_n1519), .B0(new_n1063), .Y(new_n1520));
  INV1_HPNW1   g1135(.A(new_n1071), .Y(new_n1521));
  AOI21_HPNW1  g1136(.A0(new_n1064), .A1(new_n1520), .B0(new_n1521), .Y(new_n1522));
  OAI21_HPNW1  g1137(.A0(new_n1075), .A1(new_n1522), .B0(new_n1079), .Y(new_n1523));
  INV1_HPNW1   g1138(.A(new_n1087), .Y(new_n1524));
  AOI21_HPNW1  g1139(.A0(new_n1080), .A1(new_n1523), .B0(new_n1524), .Y(new_n1525));
  OAI21_HPNW1  g1140(.A0(new_n1091), .A1(new_n1525), .B0(new_n1095), .Y(new_n1526));
  INV1_HPNW1   g1141(.A(new_n1103), .Y(new_n1527));
  AOI21_HPNW1  g1142(.A0(new_n1096), .A1(new_n1526), .B0(new_n1527), .Y(new_n1528));
  OAI21_HPNW1  g1143(.A0(new_n1107), .A1(new_n1528), .B0(new_n1111), .Y(new_n1529));
  INV1_HPNW1   g1144(.A(new_n1119), .Y(new_n1530));
  AOI21_HPNW1  g1145(.A0(new_n1112), .A1(new_n1529), .B0(new_n1530), .Y(new_n1531));
  OAI21_HPNW1  g1146(.A0(new_n1123), .A1(new_n1531), .B0(new_n1127), .Y(new_n1532));
  INV1_HPNW1   g1147(.A(new_n1135), .Y(new_n1533));
  AOI21_HPNW1  g1148(.A0(new_n1128), .A1(new_n1532), .B0(new_n1533), .Y(new_n1534));
  OAI21_HPNW1  g1149(.A0(new_n1139), .A1(new_n1534), .B0(new_n1143), .Y(new_n1535));
  INV1_HPNW1   g1150(.A(new_n1151), .Y(new_n1536));
  AOI21_HPNW1  g1151(.A0(new_n1144), .A1(new_n1535), .B0(new_n1536), .Y(new_n1537));
  OAI21_HPNW1  g1152(.A0(new_n1155), .A1(new_n1537), .B0(new_n1159), .Y(new_n1538));
  INV1_HPNW1   g1153(.A(new_n1167), .Y(new_n1539));
  AOI21_HPNW1  g1154(.A0(new_n1160), .A1(new_n1538), .B0(new_n1539), .Y(new_n1540));
  OAI21_HPNW1  g1155(.A0(new_n1171), .A1(new_n1540), .B0(new_n1175), .Y(new_n1541));
  INV1_HPNW1   g1156(.A(new_n1183), .Y(new_n1542));
  AOI21_HPNW1  g1157(.A0(new_n1176), .A1(new_n1541), .B0(new_n1542), .Y(new_n1543));
  OAI21_HPNW1  g1158(.A0(new_n1187), .A1(new_n1543), .B0(new_n1191), .Y(new_n1544));
  INV1_HPNW1   g1159(.A(new_n1199), .Y(new_n1545));
  AOI21_HPNW1  g1160(.A0(new_n1192), .A1(new_n1544), .B0(new_n1545), .Y(new_n1546));
  OAI21_HPNW1  g1161(.A0(new_n1203), .A1(new_n1546), .B0(new_n1207), .Y(new_n1547));
  INV1_HPNW1   g1162(.A(new_n1215), .Y(new_n1548));
  AOI21_HPNW1  g1163(.A0(new_n1208), .A1(new_n1547), .B0(new_n1548), .Y(new_n1549));
  OAI21_HPNW1  g1164(.A0(new_n1219), .A1(new_n1549), .B0(new_n1223), .Y(new_n1550));
  INV1_HPNW1   g1165(.A(new_n1231), .Y(new_n1551));
  AOI21_HPNW1  g1166(.A0(new_n1224), .A1(new_n1550), .B0(new_n1551), .Y(new_n1552));
  OAI21_HPNW1  g1167(.A0(new_n1235), .A1(new_n1552), .B0(new_n1239), .Y(new_n1553));
  INV1_HPNW1   g1168(.A(new_n1247), .Y(new_n1554));
  AOI21_HPNW1  g1169(.A0(new_n1240), .A1(new_n1553), .B0(new_n1554), .Y(new_n1555));
  OAI21_HPNW1  g1170(.A0(new_n1251), .A1(new_n1555), .B0(new_n1255), .Y(new_n1556));
  INV1_HPNW1   g1171(.A(new_n1263), .Y(new_n1557));
  AOI21_HPNW1  g1172(.A0(new_n1256), .A1(new_n1556), .B0(new_n1557), .Y(new_n1558));
  OAI21_HPNW1  g1173(.A0(new_n1267), .A1(new_n1558), .B0(new_n1271), .Y(new_n1559));
  INV1_HPNW1   g1174(.A(new_n1279), .Y(new_n1560));
  AOI21_HPNW1  g1175(.A0(new_n1272), .A1(new_n1559), .B0(new_n1560), .Y(new_n1561));
  OAI21_HPNW1  g1176(.A0(new_n1283), .A1(new_n1561), .B0(new_n1287), .Y(new_n1562));
  INV1_HPNW1   g1177(.A(new_n1295), .Y(new_n1563));
  AOI21_HPNW1  g1178(.A0(new_n1288), .A1(new_n1562), .B0(new_n1563), .Y(new_n1564));
  OAI21_HPNW1  g1179(.A0(new_n1299), .A1(new_n1564), .B0(new_n1303), .Y(new_n1565));
  INV1_HPNW1   g1180(.A(new_n1311), .Y(new_n1566));
  AOI21_HPNW1  g1181(.A0(new_n1304), .A1(new_n1565), .B0(new_n1566), .Y(new_n1567));
  OAI21_HPNW1  g1182(.A0(new_n1315), .A1(new_n1567), .B0(new_n1319), .Y(new_n1568));
  INV1_HPNW1   g1183(.A(new_n1327), .Y(new_n1569));
  AOI21_HPNW1  g1184(.A0(new_n1320), .A1(new_n1568), .B0(new_n1569), .Y(new_n1570));
  OAI21_HPNW1  g1185(.A0(new_n1331), .A1(new_n1570), .B0(new_n1335), .Y(new_n1571));
  INV1_HPNW1   g1186(.A(new_n1343), .Y(new_n1572));
  AOI21_HPNW1  g1187(.A0(new_n1336), .A1(new_n1571), .B0(new_n1572), .Y(new_n1573));
  OAI21_HPNW1  g1188(.A0(new_n1347), .A1(new_n1573), .B0(new_n1351), .Y(new_n1574));
  INV1_HPNW1   g1189(.A(new_n1359), .Y(new_n1575));
  AOI21_HPNW1  g1190(.A0(new_n1352), .A1(new_n1574), .B0(new_n1575), .Y(new_n1576));
  OAI21_HPNW1  g1191(.A0(new_n1363), .A1(new_n1576), .B0(new_n1367), .Y(new_n1577));
  INV1_HPNW1   g1192(.A(new_n1375), .Y(new_n1578));
  AOI21_HPNW1  g1193(.A0(new_n1368), .A1(new_n1577), .B0(new_n1578), .Y(new_n1579));
  OAI21_HPNW1  g1194(.A0(new_n1386), .A1(new_n1579), .B0(new_n1383), .Y(new_n1580));
  INV1_HPNW1   g1195(.A(new_n1393), .Y(new_n1581));
  AOI21_HPNW1  g1196(.A0(new_n1384), .A1(new_n1580), .B0(new_n1581), .Y(new_n1582));
  NOR2_HPNW1   g1197(.A(new_n1394), .B(new_n1582), .Y(\f[127] ));
  INV1_HPNW1   g1198(.A(new_n1392), .Y(new_n1584));
  NOR2_HPNW1   g1199(.A(\b[127] ), .B(\a[127] ), .Y(new_n1585));
  NAND2_HPNW1  g1200(.A(\b[127] ), .B(\a[127] ), .Y(new_n1586));
  OAI21_HPNW1  g1201(.A0(new_n1585), .A1(new_n1584), .B0(new_n1586), .Y(cOut));
endmodule


